module SimpleLACore(
  input         clock,
  input         reset,
  input         io_ipi,
  input  [7:0]  io_interrupt,
  output        io_inst_req_valid,
  output [31:0] io_inst_req_bits_addr,
  input         io_inst_resp_valid,
  input  [31:0] io_inst_resp_bits,
  output        io_data_req_valid,
  output [3:0]  io_data_req_bits_wen,
  output [31:0] io_data_req_bits_addr,
  output [31:0] io_data_req_bits_wdata,
  output        io_data_req_bits_cacop,
  output        io_data_req_bits_preld,
  input         io_data_resp_valid,
  input  [31:0] io_data_resp_bits,
  output [31:0] io_debug_pc,
  output [3:0]  io_debug_wen,
  output [4:0]  io_debug_wnum,
  output [31:0] io_debug_wdata,
  output [31:0] io_debug_inst
);
  reg [31:0] GR [0:31];
  wire  GR_rj_MPORT_en;
  wire [4:0] GR_rj_MPORT_addr;
  wire [31:0] GR_rj_MPORT_data;
  wire  GR_rkd_MPORT_en;
  wire [4:0] GR_rkd_MPORT_addr;
  wire [31:0] GR_rkd_MPORT_data;
  wire [31:0] GR_MPORT_data;
  wire [4:0] GR_MPORT_addr;
  wire  GR_MPORT_mask;
  wire  GR_MPORT_en;
  reg  idle;
  reg [31:0] PC;
  wire [31:0] PC4 = PC + 32'h4;
  reg [63:0] timer;
  wire [63:0] _timer_T_1 = timer + 64'h1;
  reg  iStallReg;
  reg  dStallReg;
  reg [1:0] crmd_DATM;
  reg [1:0] crmd_DATF;
  reg  crmd_PG;
  reg  crmd_DA;
  reg  crmd_IE;
  reg [1:0] crmd_PLV;
  reg  csrs_1_PIE;
  reg [1:0] csrs_1_PPLV;
  reg  csrs_2_FPE;
  reg [12:0] csrs_3_LIE;
  reg [5:0] csrs_4_Ecode;
  reg  csrs_4_IS_0;
  reg  csrs_4_IS_1;
  reg  csrs_4_IS_2;
  reg  csrs_4_IS_3;
  reg  csrs_4_IS_4;
  reg  csrs_4_IS_5;
  reg  csrs_4_IS_6;
  reg  csrs_4_IS_7;
  reg  csrs_4_IS_8;
  reg  csrs_4_IS_9;
  reg  csrs_4_IS_11;
  reg  csrs_4_IS_12;
  reg [31:0] csrs_5_PC;
  reg [31:0] badv_VAddr;
  reg [25:0] csrs_7_VA;
  reg  csrs_8_NE;
  reg [5:0] csrs_8_PS;
  reg [3:0] csrs_8_Index;
  reg [18:0] csrs_9_VPPN;
  reg [23:0] csrs_10_PPN;
  reg  csrs_10_G;
  reg [1:0] csrs_10_MAT;
  reg [1:0] csrs_10_PLV;
  reg  csrs_10_D;
  reg  csrs_10_V;
  reg [23:0] csrs_11_PPN;
  reg  csrs_11_G;
  reg [1:0] csrs_11_MAT;
  reg [1:0] csrs_11_PLV;
  reg  csrs_11_D;
  reg  csrs_11_V;
  reg [9:0] asid_ASID;
  reg [19:0] csrs_13_Base;
  reg [19:0] csrs_14_Base;
  reg [31:0] csrs_17_Data;
  reg [31:0] csrs_18_Data;
  reg [31:0] csrs_19_Data;
  reg [31:0] csrs_20_Data;
  reg [31:0] csrs_21_TID;
  reg [29:0] csrs_22_InitVal;
  reg  csrs_22_Periodic;
  reg  csrs_22_En;
  reg [31:0] csrs_23_TimeVal;
  reg  csrs_25_KLO;
  reg  csrs_25_ROLLB;
  reg [25:0] csrs_26_PA;
  reg [2:0] csrs_27_VSEG;
  reg [2:0] csrs_27_PSEG;
  reg [1:0] csrs_27_MAT;
  reg  csrs_27_PLV3;
  reg  csrs_27_PLV0;
  reg [2:0] csrs_28_VSEG;
  reg [2:0] csrs_28_PSEG;
  reg [1:0] csrs_28_MAT;
  reg  csrs_28_PLV3;
  reg  csrs_28_PLV0;
  wire [31:0] _tval_TimeVal_T_1 = csrs_23_TimeVal - 32'h1;
  wire  _GEN_0 = csrs_23_TimeVal == 32'h1 | csrs_4_IS_11;
  wire [31:0] _tval_TimeVal_T_2 = {csrs_22_InitVal,2'h0};
  wire [31:0] _GEN_1 = csrs_22_Periodic ? _tval_TimeVal_T_2 : csrs_23_TimeVal;
  wire [31:0] _GEN_2 = csrs_23_TimeVal != 32'h0 ? _tval_TimeVal_T_1 : _GEN_1;
  wire  _GEN_3 = csrs_23_TimeVal != 32'h0 ? _GEN_0 : csrs_4_IS_11;
  wire [31:0] _GEN_4 = csrs_22_En ? _GEN_2 : csrs_23_TimeVal;
  wire  _GEN_5 = csrs_22_En ? _GEN_3 : csrs_4_IS_11;
  wire [5:0] INT_lo = {csrs_4_IS_5,csrs_4_IS_4,csrs_4_IS_3,csrs_4_IS_2,csrs_4_IS_1,csrs_4_IS_0};
  wire [12:0] _INT_T = {csrs_4_IS_12,csrs_4_IS_11,1'h0,csrs_4_IS_9,csrs_4_IS_8,csrs_4_IS_7,csrs_4_IS_6,INT_lo};
  wire [12:0] _INT_T_1 = csrs_3_LIE & _INT_T;
  wire  INT = |_INT_T_1 & crmd_IE;
  wire  _T_28 = ~idle;
  wire  _T_31 = PC[1:0] != 2'h0;
  wire  _T_12 = crmd_PLV == 2'h0;
  wire  _T_14 = crmd_PLV == 2'h3;
  reg  tlb_0_E;
  reg [18:0] tlb_0_VPPN;
  reg [5:0] tlb_0_PS;
  wire  vaMatch_0 = tlb_0_VPPN[18:9] == PC[31:22] & (tlb_0_PS == 6'h15 | tlb_0_VPPN[8:0] == PC[21:13]);
  reg  tlb_0_G;
  reg [9:0] tlb_0_ASID;
  wire  asidMatch_0 = tlb_0_ASID == asid_ASID;
  wire  tlbHit_0 = tlb_0_E & vaMatch_0 & (tlb_0_G | asidMatch_0);
  reg  tlb_1_E;
  reg [18:0] tlb_1_VPPN;
  reg [5:0] tlb_1_PS;
  wire  vaMatch_1 = tlb_1_VPPN[18:9] == PC[31:22] & (tlb_1_PS == 6'h15 | tlb_1_VPPN[8:0] == PC[21:13]);
  reg  tlb_1_G;
  reg [9:0] tlb_1_ASID;
  wire  asidMatch_1 = tlb_1_ASID == asid_ASID;
  wire  tlbHit_1 = tlb_1_E & vaMatch_1 & (tlb_1_G | asidMatch_1);
  reg  tlb_2_E;
  reg [18:0] tlb_2_VPPN;
  reg [5:0] tlb_2_PS;
  wire  vaMatch_2 = tlb_2_VPPN[18:9] == PC[31:22] & (tlb_2_PS == 6'h15 | tlb_2_VPPN[8:0] == PC[21:13]);
  reg  tlb_2_G;
  reg [9:0] tlb_2_ASID;
  wire  asidMatch_2 = tlb_2_ASID == asid_ASID;
  wire  tlbHit_2 = tlb_2_E & vaMatch_2 & (tlb_2_G | asidMatch_2);
  reg  tlb_3_E;
  reg [18:0] tlb_3_VPPN;
  reg [5:0] tlb_3_PS;
  wire  vaMatch_3 = tlb_3_VPPN[18:9] == PC[31:22] & (tlb_3_PS == 6'h15 | tlb_3_VPPN[8:0] == PC[21:13]);
  reg  tlb_3_G;
  reg [9:0] tlb_3_ASID;
  wire  asidMatch_3 = tlb_3_ASID == asid_ASID;
  wire  tlbHit_3 = tlb_3_E & vaMatch_3 & (tlb_3_G | asidMatch_3);
  reg  tlb_4_E;
  reg [18:0] tlb_4_VPPN;
  reg [5:0] tlb_4_PS;
  wire  vaMatch_4 = tlb_4_VPPN[18:9] == PC[31:22] & (tlb_4_PS == 6'h15 | tlb_4_VPPN[8:0] == PC[21:13]);
  reg  tlb_4_G;
  reg [9:0] tlb_4_ASID;
  wire  asidMatch_4 = tlb_4_ASID == asid_ASID;
  wire  tlbHit_4 = tlb_4_E & vaMatch_4 & (tlb_4_G | asidMatch_4);
  reg  tlb_5_E;
  reg [18:0] tlb_5_VPPN;
  reg [5:0] tlb_5_PS;
  wire  vaMatch_5 = tlb_5_VPPN[18:9] == PC[31:22] & (tlb_5_PS == 6'h15 | tlb_5_VPPN[8:0] == PC[21:13]);
  reg  tlb_5_G;
  reg [9:0] tlb_5_ASID;
  wire  asidMatch_5 = tlb_5_ASID == asid_ASID;
  wire  tlbHit_5 = tlb_5_E & vaMatch_5 & (tlb_5_G | asidMatch_5);
  reg  tlb_6_E;
  reg [18:0] tlb_6_VPPN;
  reg [5:0] tlb_6_PS;
  wire  vaMatch_6 = tlb_6_VPPN[18:9] == PC[31:22] & (tlb_6_PS == 6'h15 | tlb_6_VPPN[8:0] == PC[21:13]);
  reg  tlb_6_G;
  reg [9:0] tlb_6_ASID;
  wire  asidMatch_6 = tlb_6_ASID == asid_ASID;
  wire  tlbHit_6 = tlb_6_E & vaMatch_6 & (tlb_6_G | asidMatch_6);
  reg  tlb_7_E;
  reg [18:0] tlb_7_VPPN;
  reg [5:0] tlb_7_PS;
  wire  vaMatch_7 = tlb_7_VPPN[18:9] == PC[31:22] & (tlb_7_PS == 6'h15 | tlb_7_VPPN[8:0] == PC[21:13]);
  reg  tlb_7_G;
  reg [9:0] tlb_7_ASID;
  wire  asidMatch_7 = tlb_7_ASID == asid_ASID;
  wire  tlbHit_7 = tlb_7_E & vaMatch_7 & (tlb_7_G | asidMatch_7);
  reg  tlb_8_E;
  reg [18:0] tlb_8_VPPN;
  reg [5:0] tlb_8_PS;
  wire  vaMatch_8 = tlb_8_VPPN[18:9] == PC[31:22] & (tlb_8_PS == 6'h15 | tlb_8_VPPN[8:0] == PC[21:13]);
  reg  tlb_8_G;
  reg [9:0] tlb_8_ASID;
  wire  asidMatch_8 = tlb_8_ASID == asid_ASID;
  wire  tlbHit_8 = tlb_8_E & vaMatch_8 & (tlb_8_G | asidMatch_8);
  reg  tlb_9_E;
  reg [18:0] tlb_9_VPPN;
  reg [5:0] tlb_9_PS;
  wire  vaMatch_9 = tlb_9_VPPN[18:9] == PC[31:22] & (tlb_9_PS == 6'h15 | tlb_9_VPPN[8:0] == PC[21:13]);
  reg  tlb_9_G;
  reg [9:0] tlb_9_ASID;
  wire  asidMatch_9 = tlb_9_ASID == asid_ASID;
  wire  tlbHit_9 = tlb_9_E & vaMatch_9 & (tlb_9_G | asidMatch_9);
  reg  tlb_10_E;
  reg [18:0] tlb_10_VPPN;
  reg [5:0] tlb_10_PS;
  wire  vaMatch_10 = tlb_10_VPPN[18:9] == PC[31:22] & (tlb_10_PS == 6'h15 | tlb_10_VPPN[8:0] == PC[21:13]);
  reg  tlb_10_G;
  reg [9:0] tlb_10_ASID;
  wire  asidMatch_10 = tlb_10_ASID == asid_ASID;
  wire  tlbHit_10 = tlb_10_E & vaMatch_10 & (tlb_10_G | asidMatch_10);
  reg  tlb_11_E;
  reg [18:0] tlb_11_VPPN;
  reg [5:0] tlb_11_PS;
  wire  vaMatch_11 = tlb_11_VPPN[18:9] == PC[31:22] & (tlb_11_PS == 6'h15 | tlb_11_VPPN[8:0] == PC[21:13]);
  reg  tlb_11_G;
  reg [9:0] tlb_11_ASID;
  wire  asidMatch_11 = tlb_11_ASID == asid_ASID;
  wire  tlbHit_11 = tlb_11_E & vaMatch_11 & (tlb_11_G | asidMatch_11);
  reg  tlb_12_E;
  reg [18:0] tlb_12_VPPN;
  reg [5:0] tlb_12_PS;
  wire  vaMatch_12 = tlb_12_VPPN[18:9] == PC[31:22] & (tlb_12_PS == 6'h15 | tlb_12_VPPN[8:0] == PC[21:13]);
  reg  tlb_12_G;
  reg [9:0] tlb_12_ASID;
  wire  asidMatch_12 = tlb_12_ASID == asid_ASID;
  wire  tlbHit_12 = tlb_12_E & vaMatch_12 & (tlb_12_G | asidMatch_12);
  reg  tlb_13_E;
  reg [18:0] tlb_13_VPPN;
  reg [5:0] tlb_13_PS;
  wire  vaMatch_13 = tlb_13_VPPN[18:9] == PC[31:22] & (tlb_13_PS == 6'h15 | tlb_13_VPPN[8:0] == PC[21:13]);
  reg  tlb_13_G;
  reg [9:0] tlb_13_ASID;
  wire  asidMatch_13 = tlb_13_ASID == asid_ASID;
  wire  tlbHit_13 = tlb_13_E & vaMatch_13 & (tlb_13_G | asidMatch_13);
  reg  tlb_14_E;
  reg [18:0] tlb_14_VPPN;
  reg [5:0] tlb_14_PS;
  wire  vaMatch_14 = tlb_14_VPPN[18:9] == PC[31:22] & (tlb_14_PS == 6'h15 | tlb_14_VPPN[8:0] == PC[21:13]);
  reg  tlb_14_G;
  reg [9:0] tlb_14_ASID;
  wire  asidMatch_14 = tlb_14_ASID == asid_ASID;
  wire  tlbHit_14 = tlb_14_E & vaMatch_14 & (tlb_14_G | asidMatch_14);
  reg  tlb_15_E;
  reg [18:0] tlb_15_VPPN;
  reg [5:0] tlb_15_PS;
  wire  vaMatch_15 = tlb_15_VPPN[18:9] == PC[31:22] & (tlb_15_PS == 6'h15 | tlb_15_VPPN[8:0] == PC[21:13]);
  reg  tlb_15_G;
  reg [9:0] tlb_15_ASID;
  wire  asidMatch_15 = tlb_15_ASID == asid_ASID;
  wire  tlbHit_15 = tlb_15_E & vaMatch_15 & (tlb_15_G | asidMatch_15);
  wire  _GEN_9 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : ~(tlbHit_0 |
    tlbHit_1 | tlbHit_2 | tlbHit_3 | tlbHit_4 | tlbHit_5 | tlbHit_6 | tlbHit_7 | tlbHit_8 | tlbHit_9 | tlbHit_10 |
    tlbHit_11 | tlbHit_12 | tlbHit_13 | tlbHit_14 | tlbHit_15);
  wire  miss = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0 :
    _GEN_9;
  wire  _GEN_36 = crmd_DA ? 1'h0 : miss;
  wire  _GEN_41 = PC[1:0] != 2'h0 ? 1'h0 : _GEN_36;
  wire  _GEN_49 = ~INT & ~idle & _GEN_41;
  wire  _GEN_56 = dStallReg | iStallReg ? 1'h0 : _GEN_49;
  wire [5:0] _foundTLB_T_403 = tlbHit_0 ? tlb_0_PS : 6'h0;
  wire [5:0] _foundTLB_T_404 = tlbHit_1 ? tlb_1_PS : 6'h0;
  wire [5:0] _foundTLB_T_419 = _foundTLB_T_403 | _foundTLB_T_404;
  wire [5:0] _foundTLB_T_405 = tlbHit_2 ? tlb_2_PS : 6'h0;
  wire [5:0] _foundTLB_T_420 = _foundTLB_T_419 | _foundTLB_T_405;
  wire [5:0] _foundTLB_T_406 = tlbHit_3 ? tlb_3_PS : 6'h0;
  wire [5:0] _foundTLB_T_421 = _foundTLB_T_420 | _foundTLB_T_406;
  wire [5:0] _foundTLB_T_407 = tlbHit_4 ? tlb_4_PS : 6'h0;
  wire [5:0] _foundTLB_T_422 = _foundTLB_T_421 | _foundTLB_T_407;
  wire [5:0] _foundTLB_T_408 = tlbHit_5 ? tlb_5_PS : 6'h0;
  wire [5:0] _foundTLB_T_423 = _foundTLB_T_422 | _foundTLB_T_408;
  wire [5:0] _foundTLB_T_409 = tlbHit_6 ? tlb_6_PS : 6'h0;
  wire [5:0] _foundTLB_T_424 = _foundTLB_T_423 | _foundTLB_T_409;
  wire [5:0] _foundTLB_T_410 = tlbHit_7 ? tlb_7_PS : 6'h0;
  wire [5:0] _foundTLB_T_425 = _foundTLB_T_424 | _foundTLB_T_410;
  wire [5:0] _foundTLB_T_411 = tlbHit_8 ? tlb_8_PS : 6'h0;
  wire [5:0] _foundTLB_T_426 = _foundTLB_T_425 | _foundTLB_T_411;
  wire [5:0] _foundTLB_T_412 = tlbHit_9 ? tlb_9_PS : 6'h0;
  wire [5:0] _foundTLB_T_427 = _foundTLB_T_426 | _foundTLB_T_412;
  wire [5:0] _foundTLB_T_413 = tlbHit_10 ? tlb_10_PS : 6'h0;
  wire [5:0] _foundTLB_T_428 = _foundTLB_T_427 | _foundTLB_T_413;
  wire [5:0] _foundTLB_T_414 = tlbHit_11 ? tlb_11_PS : 6'h0;
  wire [5:0] _foundTLB_T_429 = _foundTLB_T_428 | _foundTLB_T_414;
  wire [5:0] _foundTLB_T_415 = tlbHit_12 ? tlb_12_PS : 6'h0;
  wire [5:0] _foundTLB_T_430 = _foundTLB_T_429 | _foundTLB_T_415;
  wire [5:0] _foundTLB_T_416 = tlbHit_13 ? tlb_13_PS : 6'h0;
  wire [5:0] _foundTLB_T_431 = _foundTLB_T_430 | _foundTLB_T_416;
  wire [5:0] _foundTLB_T_417 = tlbHit_14 ? tlb_14_PS : 6'h0;
  wire [5:0] _foundTLB_T_432 = _foundTLB_T_431 | _foundTLB_T_417;
  wire [5:0] _foundTLB_T_418 = tlbHit_15 ? tlb_15_PS : 6'h0;
  wire [5:0] foundTLB_PS = _foundTLB_T_432 | _foundTLB_T_418;
  wire  _oddPG_T = foundTLB_PS == 6'hc;
  wire  oddPG = foundTLB_PS == 6'hc ? PC[12] : PC[21];
  reg  tlb_0_P1_V;
  reg  tlb_1_P1_V;
  reg  tlb_2_P1_V;
  reg  tlb_3_P1_V;
  reg  tlb_4_P1_V;
  reg  tlb_5_P1_V;
  reg  tlb_6_P1_V;
  reg  tlb_7_P1_V;
  reg  tlb_8_P1_V;
  reg  tlb_9_P1_V;
  reg  tlb_10_P1_V;
  reg  tlb_11_P1_V;
  reg  tlb_12_P1_V;
  reg  tlb_13_P1_V;
  reg  tlb_14_P1_V;
  reg  tlb_15_P1_V;
  wire  _foundTLB_T_15 = tlbHit_15 & tlb_15_P1_V;
  wire  foundTLB_P1_V = tlbHit_0 & tlb_0_P1_V | tlbHit_1 & tlb_1_P1_V | tlbHit_2 & tlb_2_P1_V | tlbHit_3 & tlb_3_P1_V |
    tlbHit_4 & tlb_4_P1_V | tlbHit_5 & tlb_5_P1_V | tlbHit_6 & tlb_6_P1_V | tlbHit_7 & tlb_7_P1_V | tlbHit_8 &
    tlb_8_P1_V | tlbHit_9 & tlb_9_P1_V | tlbHit_10 & tlb_10_P1_V | tlbHit_11 & tlb_11_P1_V | tlbHit_12 & tlb_12_P1_V |
    tlbHit_13 & tlb_13_P1_V | tlbHit_14 & tlb_14_P1_V | _foundTLB_T_15;
  reg  tlb_0_P0_V;
  reg  tlb_1_P0_V;
  reg  tlb_2_P0_V;
  reg  tlb_3_P0_V;
  reg  tlb_4_P0_V;
  reg  tlb_5_P0_V;
  reg  tlb_6_P0_V;
  reg  tlb_7_P0_V;
  reg  tlb_8_P0_V;
  reg  tlb_9_P0_V;
  reg  tlb_10_P0_V;
  reg  tlb_11_P0_V;
  reg  tlb_12_P0_V;
  reg  tlb_13_P0_V;
  reg  tlb_14_P0_V;
  reg  tlb_15_P0_V;
  wire  _foundTLB_T_170 = tlbHit_15 & tlb_15_P0_V;
  wire  foundTLB_P0_V = tlbHit_0 & tlb_0_P0_V | tlbHit_1 & tlb_1_P0_V | tlbHit_2 & tlb_2_P0_V | tlbHit_3 & tlb_3_P0_V |
    tlbHit_4 & tlb_4_P0_V | tlbHit_5 & tlb_5_P0_V | tlbHit_6 & tlb_6_P0_V | tlbHit_7 & tlb_7_P0_V | tlbHit_8 &
    tlb_8_P0_V | tlbHit_9 & tlb_9_P0_V | tlbHit_10 & tlb_10_P0_V | tlbHit_11 & tlb_11_P0_V | tlbHit_12 & tlb_12_P0_V |
    tlbHit_13 & tlb_13_P0_V | tlbHit_14 & tlb_14_P0_V | _foundTLB_T_170;
  wire  foundP_V = oddPG ? foundTLB_P1_V : foundTLB_P0_V;
  wire  _GEN_10 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : ~foundP_V;
  wire  invalid = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_10;
  reg [1:0] tlb_0_P1_PLV;
  wire [1:0] _foundTLB_T_93 = tlbHit_0 ? tlb_0_P1_PLV : 2'h0;
  reg [1:0] tlb_1_P1_PLV;
  wire [1:0] _foundTLB_T_94 = tlbHit_1 ? tlb_1_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_109 = _foundTLB_T_93 | _foundTLB_T_94;
  reg [1:0] tlb_2_P1_PLV;
  wire [1:0] _foundTLB_T_95 = tlbHit_2 ? tlb_2_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_110 = _foundTLB_T_109 | _foundTLB_T_95;
  reg [1:0] tlb_3_P1_PLV;
  wire [1:0] _foundTLB_T_96 = tlbHit_3 ? tlb_3_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_111 = _foundTLB_T_110 | _foundTLB_T_96;
  reg [1:0] tlb_4_P1_PLV;
  wire [1:0] _foundTLB_T_97 = tlbHit_4 ? tlb_4_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_112 = _foundTLB_T_111 | _foundTLB_T_97;
  reg [1:0] tlb_5_P1_PLV;
  wire [1:0] _foundTLB_T_98 = tlbHit_5 ? tlb_5_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_113 = _foundTLB_T_112 | _foundTLB_T_98;
  reg [1:0] tlb_6_P1_PLV;
  wire [1:0] _foundTLB_T_99 = tlbHit_6 ? tlb_6_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_114 = _foundTLB_T_113 | _foundTLB_T_99;
  reg [1:0] tlb_7_P1_PLV;
  wire [1:0] _foundTLB_T_100 = tlbHit_7 ? tlb_7_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_115 = _foundTLB_T_114 | _foundTLB_T_100;
  reg [1:0] tlb_8_P1_PLV;
  wire [1:0] _foundTLB_T_101 = tlbHit_8 ? tlb_8_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_116 = _foundTLB_T_115 | _foundTLB_T_101;
  reg [1:0] tlb_9_P1_PLV;
  wire [1:0] _foundTLB_T_102 = tlbHit_9 ? tlb_9_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_117 = _foundTLB_T_116 | _foundTLB_T_102;
  reg [1:0] tlb_10_P1_PLV;
  wire [1:0] _foundTLB_T_103 = tlbHit_10 ? tlb_10_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_118 = _foundTLB_T_117 | _foundTLB_T_103;
  reg [1:0] tlb_11_P1_PLV;
  wire [1:0] _foundTLB_T_104 = tlbHit_11 ? tlb_11_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_119 = _foundTLB_T_118 | _foundTLB_T_104;
  reg [1:0] tlb_12_P1_PLV;
  wire [1:0] _foundTLB_T_105 = tlbHit_12 ? tlb_12_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_120 = _foundTLB_T_119 | _foundTLB_T_105;
  reg [1:0] tlb_13_P1_PLV;
  wire [1:0] _foundTLB_T_106 = tlbHit_13 ? tlb_13_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_121 = _foundTLB_T_120 | _foundTLB_T_106;
  reg [1:0] tlb_14_P1_PLV;
  wire [1:0] _foundTLB_T_107 = tlbHit_14 ? tlb_14_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_122 = _foundTLB_T_121 | _foundTLB_T_107;
  reg [1:0] tlb_15_P1_PLV;
  wire [1:0] _foundTLB_T_108 = tlbHit_15 ? tlb_15_P1_PLV : 2'h0;
  wire [1:0] foundTLB_P1_PLV = _foundTLB_T_122 | _foundTLB_T_108;
  reg [1:0] tlb_0_P0_PLV;
  wire [1:0] _foundTLB_T_248 = tlbHit_0 ? tlb_0_P0_PLV : 2'h0;
  reg [1:0] tlb_1_P0_PLV;
  wire [1:0] _foundTLB_T_249 = tlbHit_1 ? tlb_1_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_264 = _foundTLB_T_248 | _foundTLB_T_249;
  reg [1:0] tlb_2_P0_PLV;
  wire [1:0] _foundTLB_T_250 = tlbHit_2 ? tlb_2_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_265 = _foundTLB_T_264 | _foundTLB_T_250;
  reg [1:0] tlb_3_P0_PLV;
  wire [1:0] _foundTLB_T_251 = tlbHit_3 ? tlb_3_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_266 = _foundTLB_T_265 | _foundTLB_T_251;
  reg [1:0] tlb_4_P0_PLV;
  wire [1:0] _foundTLB_T_252 = tlbHit_4 ? tlb_4_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_267 = _foundTLB_T_266 | _foundTLB_T_252;
  reg [1:0] tlb_5_P0_PLV;
  wire [1:0] _foundTLB_T_253 = tlbHit_5 ? tlb_5_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_268 = _foundTLB_T_267 | _foundTLB_T_253;
  reg [1:0] tlb_6_P0_PLV;
  wire [1:0] _foundTLB_T_254 = tlbHit_6 ? tlb_6_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_269 = _foundTLB_T_268 | _foundTLB_T_254;
  reg [1:0] tlb_7_P0_PLV;
  wire [1:0] _foundTLB_T_255 = tlbHit_7 ? tlb_7_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_270 = _foundTLB_T_269 | _foundTLB_T_255;
  reg [1:0] tlb_8_P0_PLV;
  wire [1:0] _foundTLB_T_256 = tlbHit_8 ? tlb_8_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_271 = _foundTLB_T_270 | _foundTLB_T_256;
  reg [1:0] tlb_9_P0_PLV;
  wire [1:0] _foundTLB_T_257 = tlbHit_9 ? tlb_9_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_272 = _foundTLB_T_271 | _foundTLB_T_257;
  reg [1:0] tlb_10_P0_PLV;
  wire [1:0] _foundTLB_T_258 = tlbHit_10 ? tlb_10_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_273 = _foundTLB_T_272 | _foundTLB_T_258;
  reg [1:0] tlb_11_P0_PLV;
  wire [1:0] _foundTLB_T_259 = tlbHit_11 ? tlb_11_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_274 = _foundTLB_T_273 | _foundTLB_T_259;
  reg [1:0] tlb_12_P0_PLV;
  wire [1:0] _foundTLB_T_260 = tlbHit_12 ? tlb_12_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_275 = _foundTLB_T_274 | _foundTLB_T_260;
  reg [1:0] tlb_13_P0_PLV;
  wire [1:0] _foundTLB_T_261 = tlbHit_13 ? tlb_13_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_276 = _foundTLB_T_275 | _foundTLB_T_261;
  reg [1:0] tlb_14_P0_PLV;
  wire [1:0] _foundTLB_T_262 = tlbHit_14 ? tlb_14_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_277 = _foundTLB_T_276 | _foundTLB_T_262;
  reg [1:0] tlb_15_P0_PLV;
  wire [1:0] _foundTLB_T_263 = tlbHit_15 ? tlb_15_P0_PLV : 2'h0;
  wire [1:0] foundTLB_P0_PLV = _foundTLB_T_277 | _foundTLB_T_263;
  wire [1:0] foundP_PLV = oddPG ? foundTLB_P1_PLV : foundTLB_P0_PLV;
  wire  _GEN_11 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : crmd_PLV >
    foundP_PLV;
  wire  ppi = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0 :
    _GEN_11;
  wire  _GEN_21 = ppi ? 1'h0 : 1'h1;
  wire  _GEN_24 = invalid ? 1'h0 : _GEN_21;
  wire  _GEN_28 = miss ? 1'h0 : _GEN_24;
  wire  _GEN_34 = crmd_DA | _GEN_28;
  wire  _GEN_40 = PC[1:0] != 2'h0 ? 1'h0 : _GEN_34;
  wire  _GEN_48 = ~INT & ~idle & _GEN_40;
  wire  IF_OK = dStallReg | iStallReg | _GEN_48;
  wire  iStall = ~io_inst_resp_valid & (io_inst_req_valid | iStallReg);
  wire  _T_1316 = ~iStall;
  reg [31:0] inst_reg;
  wire [31:0] inst = dStallReg ? inst_reg : io_inst_resp_bits;
  wire [31:0] _T_34 = inst & 32'hfffffc1f;
  wire  _T_35 = 32'h6000 == _T_34;
  wire [31:0] _T_36 = inst & 32'hffffffe0;
  wire  _T_37 = 32'h6000 == _T_36;
  wire  _T_39 = 32'h6400 == _T_36;
  wire [31:0] _T_40 = inst & 32'hffff8000;
  wire  _T_41 = 32'h100000 == _T_40;
  wire  _T_43 = 32'h110000 == _T_40;
  wire  _T_45 = 32'h120000 == _T_40;
  wire  _T_47 = 32'h128000 == _T_40;
  wire  _T_49 = 32'h140000 == _T_40;
  wire  _T_51 = 32'h148000 == _T_40;
  wire  _T_53 = 32'h150000 == _T_40;
  wire  _T_55 = 32'h158000 == _T_40;
  wire  _T_57 = 32'h170000 == _T_40;
  wire  _T_59 = 32'h178000 == _T_40;
  wire  _T_61 = 32'h180000 == _T_40;
  wire  _T_63 = 32'h1c0000 == _T_40;
  wire  _T_65 = 32'h1c8000 == _T_40;
  wire  _T_67 = 32'h1d0000 == _T_40;
  wire  _T_69 = 32'h200000 == _T_40;
  wire  _T_71 = 32'h208000 == _T_40;
  wire  _T_73 = 32'h210000 == _T_40;
  wire  _T_75 = 32'h218000 == _T_40;
  wire  _T_77 = 32'h2a0000 == _T_40;
  wire  _T_79 = 32'h2b0000 == _T_40;
  wire  _T_81 = 32'h408000 == _T_40;
  wire  _T_83 = 32'h448000 == _T_40;
  wire  _T_85 = 32'h488000 == _T_40;
  wire [31:0] _T_86 = inst & 32'hffc00000;
  wire  _T_87 = 32'h2000000 == _T_86;
  wire  _T_89 = 32'h2400000 == _T_86;
  wire  _T_91 = 32'h2800000 == _T_86;
  wire  _T_93 = 32'h3400000 == _T_86;
  wire  _T_95 = 32'h3800000 == _T_86;
  wire  _T_97 = 32'h3c00000 == _T_86;
  wire [31:0] _T_98 = inst & 32'hff000000;
  wire  _T_99 = 32'h4000000 == _T_98;
  wire  _T_101 = 32'h6000000 == _T_86;
  wire  _T_103 = 32'h6482800 == inst;
  wire  _T_105 = 32'h6482c00 == inst;
  wire  _T_107 = 32'h6483000 == inst;
  wire  _T_109 = 32'h6483400 == inst;
  wire  _T_111 = 32'h6498000 == _T_40;
  wire  _T_113 = 32'h6483800 == inst;
  wire  _T_115 = 32'h6488000 == _T_40;
  wire [31:0] _T_116 = inst & 32'hfe000000;
  wire  _T_117 = 32'h14000000 == _T_116;
  wire  _T_119 = 32'h1c000000 == _T_116;
  wire  _T_121 = 32'h20000000 == _T_98;
  wire  _T_123 = 32'h21000000 == _T_98;
  wire  _T_125 = 32'h28000000 == _T_86;
  wire  _T_127 = 32'h28400000 == _T_86;
  wire  _T_129 = 32'h28800000 == _T_86;
  wire  _T_131 = 32'h29000000 == _T_86;
  wire  _T_133 = 32'h29400000 == _T_86;
  wire  _T_135 = 32'h29800000 == _T_86;
  wire  _T_137 = 32'h2a000000 == _T_86;
  wire  _T_139 = 32'h2a400000 == _T_86;
  wire  _T_141 = 32'h2ac00000 == _T_86;
  wire  _T_143 = 32'h38720000 == _T_40;
  wire  _T_145 = 32'h38728000 == _T_40;
  wire [31:0] _T_146 = inst & 32'hfc000000;
  wire  _T_147 = 32'h4c000000 == _T_146;
  wire  _T_149 = 32'h50000000 == _T_146;
  wire  _T_151 = 32'h54000000 == _T_146;
  wire  _T_153 = 32'h58000000 == _T_146;
  wire  _T_155 = 32'h5c000000 == _T_146;
  wire  _T_157 = 32'h60000000 == _T_146;
  wire  _T_159 = 32'h64000000 == _T_146;
  wire  _T_161 = 32'h68000000 == _T_146;
  wire  _T_163 = 32'h6c000000 == _T_146;
  wire  _T_911 = _T_77 ? 1'h0 : _T_79;
  wire  _T_912 = _T_75 ? 1'h0 : _T_911;
  wire  _T_913 = _T_73 ? 1'h0 : _T_912;
  wire  _T_914 = _T_71 ? 1'h0 : _T_913;
  wire  _T_915 = _T_69 ? 1'h0 : _T_914;
  wire  _T_916 = _T_67 ? 1'h0 : _T_915;
  wire  _T_917 = _T_65 ? 1'h0 : _T_916;
  wire  _T_918 = _T_63 ? 1'h0 : _T_917;
  wire  _T_919 = _T_61 ? 1'h0 : _T_918;
  wire  _T_920 = _T_59 ? 1'h0 : _T_919;
  wire  _T_921 = _T_57 ? 1'h0 : _T_920;
  wire  _T_922 = _T_55 ? 1'h0 : _T_921;
  wire  _T_923 = _T_53 ? 1'h0 : _T_922;
  wire  _T_924 = _T_51 ? 1'h0 : _T_923;
  wire  _T_925 = _T_49 ? 1'h0 : _T_924;
  wire  _T_926 = _T_47 ? 1'h0 : _T_925;
  wire  _T_927 = _T_45 ? 1'h0 : _T_926;
  wire  _T_928 = _T_43 ? 1'h0 : _T_927;
  wire  _T_929 = _T_41 ? 1'h0 : _T_928;
  wire  _T_930 = _T_39 ? 1'h0 : _T_929;
  wire  _T_931 = _T_37 ? 1'h0 : _T_930;
  wire  c0_6 = _T_35 ? 1'h0 : _T_931;
  wire  _GEN_62 = IF_OK & ~iStall & c0_6;
  wire  SYS = dStallReg ? 1'h0 : _GEN_62;
  wire  _T_848 = _T_75 ? 1'h0 : _T_77;
  wire  _T_849 = _T_73 ? 1'h0 : _T_848;
  wire  _T_850 = _T_71 ? 1'h0 : _T_849;
  wire  _T_851 = _T_69 ? 1'h0 : _T_850;
  wire  _T_852 = _T_67 ? 1'h0 : _T_851;
  wire  _T_853 = _T_65 ? 1'h0 : _T_852;
  wire  _T_854 = _T_63 ? 1'h0 : _T_853;
  wire  _T_855 = _T_61 ? 1'h0 : _T_854;
  wire  _T_856 = _T_59 ? 1'h0 : _T_855;
  wire  _T_857 = _T_57 ? 1'h0 : _T_856;
  wire  _T_858 = _T_55 ? 1'h0 : _T_857;
  wire  _T_859 = _T_53 ? 1'h0 : _T_858;
  wire  _T_860 = _T_51 ? 1'h0 : _T_859;
  wire  _T_861 = _T_49 ? 1'h0 : _T_860;
  wire  _T_862 = _T_47 ? 1'h0 : _T_861;
  wire  _T_863 = _T_45 ? 1'h0 : _T_862;
  wire  _T_864 = _T_43 ? 1'h0 : _T_863;
  wire  _T_865 = _T_41 ? 1'h0 : _T_864;
  wire  _T_866 = _T_39 ? 1'h0 : _T_865;
  wire  _T_867 = _T_37 ? 1'h0 : _T_866;
  wire  break_ = _T_35 ? 1'h0 : _T_867;
  wire  _GEN_63 = IF_OK & ~iStall & break_;
  wire  BRK = dStallReg ? 1'h0 : _GEN_63;
  wire  _T_194 = _T_103 | (_T_105 | (_T_107 | (_T_109 | (_T_111 | (_T_113 | (_T_115 | (_T_117 | (_T_119 | (_T_121 | (
    _T_123 | (_T_125 | (_T_127 | (_T_129 | (_T_131 | (_T_133 | (_T_135 | (_T_137 | (_T_139 | (_T_141 | (_T_143 | (_T_145
     | (_T_147 | (_T_149 | (_T_151 | (_T_153 | (_T_155 | (_T_157 | (_T_159 | (_T_161 | _T_163)))))))))))))))))))))))))))
    ));
  wire  _T_224 = _T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53 | (_T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (
    _T_65 | (_T_67 | (_T_69 | (_T_71 | (_T_73 | (_T_75 | (_T_77 | (_T_79 | (_T_81 | (_T_83 | (_T_85 | (_T_87 | (_T_89 |
    (_T_91 | (_T_93 | (_T_95 | (_T_97 | (_T_99 | (_T_101 | _T_194)))))))))))))))))))))))))))));
  wire  instV = _T_35 | (_T_37 | (_T_39 | (_T_41 | _T_224)));
  wire [2:0] _T_958 = _T_111 ? 3'h5 : 3'h0;
  wire [2:0] _T_959 = _T_109 ? 3'h4 : _T_958;
  wire [2:0] _T_960 = _T_107 ? 3'h3 : _T_959;
  wire [2:0] _T_961 = _T_105 ? 3'h2 : _T_960;
  wire [2:0] _T_962 = _T_103 ? 3'h1 : _T_961;
  wire [2:0] _T_963 = _T_101 ? 3'h0 : _T_962;
  wire [2:0] _T_964 = _T_99 ? 3'h0 : _T_963;
  wire [2:0] _T_965 = _T_97 ? 3'h0 : _T_964;
  wire [2:0] _T_966 = _T_95 ? 3'h0 : _T_965;
  wire [2:0] _T_967 = _T_93 ? 3'h0 : _T_966;
  wire [2:0] _T_968 = _T_91 ? 3'h0 : _T_967;
  wire [2:0] _T_969 = _T_89 ? 3'h0 : _T_968;
  wire [2:0] _T_970 = _T_87 ? 3'h0 : _T_969;
  wire [2:0] _T_971 = _T_85 ? 3'h0 : _T_970;
  wire [2:0] _T_972 = _T_83 ? 3'h0 : _T_971;
  wire [2:0] _T_973 = _T_81 ? 3'h0 : _T_972;
  wire [2:0] _T_974 = _T_79 ? 3'h0 : _T_973;
  wire [2:0] _T_975 = _T_77 ? 3'h0 : _T_974;
  wire [2:0] _T_976 = _T_75 ? 3'h0 : _T_975;
  wire [2:0] _T_977 = _T_73 ? 3'h0 : _T_976;
  wire [2:0] _T_978 = _T_71 ? 3'h0 : _T_977;
  wire [2:0] _T_979 = _T_69 ? 3'h0 : _T_978;
  wire [2:0] _T_980 = _T_67 ? 3'h0 : _T_979;
  wire [2:0] _T_981 = _T_65 ? 3'h0 : _T_980;
  wire [2:0] _T_982 = _T_63 ? 3'h0 : _T_981;
  wire [2:0] _T_983 = _T_61 ? 3'h0 : _T_982;
  wire [2:0] _T_984 = _T_59 ? 3'h0 : _T_983;
  wire [2:0] _T_985 = _T_57 ? 3'h0 : _T_984;
  wire [2:0] _T_986 = _T_55 ? 3'h0 : _T_985;
  wire [2:0] _T_987 = _T_53 ? 3'h0 : _T_986;
  wire [2:0] _T_988 = _T_51 ? 3'h0 : _T_987;
  wire [2:0] _T_989 = _T_49 ? 3'h0 : _T_988;
  wire [2:0] _T_990 = _T_47 ? 3'h0 : _T_989;
  wire [2:0] _T_991 = _T_45 ? 3'h0 : _T_990;
  wire [2:0] _T_992 = _T_43 ? 3'h0 : _T_991;
  wire [2:0] _T_993 = _T_41 ? 3'h0 : _T_992;
  wire [2:0] _T_994 = _T_39 ? 3'h0 : _T_993;
  wire [2:0] _T_995 = _T_37 ? 3'h0 : _T_994;
  wire [2:0] c0_7 = _T_35 ? 3'h0 : _T_995;
  wire  _INE_T_1 = c0_7 == 3'h5;
  wire [4:0] d = inst[4:0];
  wire  inv_op_decode_0 = d == 5'h0 | d == 5'h1;
  wire  inv_op_decode_1 = d == 5'h2;
  wire  inv_op_decode_2 = d == 5'h3;
  wire  inv_op_decode_3 = d == 5'h4;
  wire  inv_op_decode_4 = d == 5'h5;
  wire  inv_op_decode_5 = d == 5'h6;
  wire  _GEN_64 = IF_OK & ~iStall & (~instV | c0_7 == 3'h5 & ~(inv_op_decode_0 | inv_op_decode_1 | inv_op_decode_2 |
    inv_op_decode_3 | inv_op_decode_4 | inv_op_decode_5));
  wire  INE = dStallReg ? 1'h0 : _GEN_64;
  wire  _T_1322 = ~SYS & ~BRK & ~INE;
  wire  _GEN_65 = IF_OK & ~iStall & _T_1322;
  wire  ID_OK = dStallReg | _GEN_65;
  wire [2:0] _T_687 = _T_141 ? 3'h0 : 3'h7;
  wire [2:0] _T_688 = _T_139 ? 3'h3 : _T_687;
  wire [2:0] _T_689 = _T_137 ? 3'h1 : _T_688;
  wire [2:0] _T_690 = _T_135 ? 3'h4 : _T_689;
  wire [2:0] _T_691 = _T_133 ? 3'h2 : _T_690;
  wire [2:0] _T_692 = _T_131 ? 3'h0 : _T_691;
  wire [2:0] _T_693 = _T_129 ? 3'h4 : _T_692;
  wire [2:0] _T_694 = _T_127 ? 3'h2 : _T_693;
  wire [2:0] _T_695 = _T_125 ? 3'h0 : _T_694;
  wire [2:0] _T_696 = _T_123 ? 3'h4 : _T_695;
  wire [2:0] _T_697 = _T_121 ? 3'h4 : _T_696;
  wire [2:0] _T_698 = _T_119 ? 3'h7 : _T_697;
  wire [2:0] _T_699 = _T_117 ? 3'h7 : _T_698;
  wire [2:0] _T_700 = _T_115 ? 3'h7 : _T_699;
  wire [2:0] _T_701 = _T_113 ? 3'h7 : _T_700;
  wire [2:0] _T_702 = _T_111 ? 3'h7 : _T_701;
  wire [2:0] _T_703 = _T_109 ? 3'h7 : _T_702;
  wire [2:0] _T_704 = _T_107 ? 3'h7 : _T_703;
  wire [2:0] _T_705 = _T_105 ? 3'h7 : _T_704;
  wire [2:0] _T_706 = _T_103 ? 3'h7 : _T_705;
  wire [2:0] _T_707 = _T_101 ? 3'h0 : _T_706;
  wire [2:0] _T_708 = _T_99 ? 3'h7 : _T_707;
  wire [2:0] _T_709 = _T_97 ? 3'h7 : _T_708;
  wire [2:0] _T_710 = _T_95 ? 3'h7 : _T_709;
  wire [2:0] _T_711 = _T_93 ? 3'h7 : _T_710;
  wire [2:0] _T_712 = _T_91 ? 3'h7 : _T_711;
  wire [2:0] _T_713 = _T_89 ? 3'h7 : _T_712;
  wire [2:0] _T_714 = _T_87 ? 3'h7 : _T_713;
  wire [2:0] _T_715 = _T_85 ? 3'h7 : _T_714;
  wire [2:0] _T_716 = _T_83 ? 3'h7 : _T_715;
  wire [2:0] _T_717 = _T_81 ? 3'h7 : _T_716;
  wire [2:0] _T_718 = _T_79 ? 3'h7 : _T_717;
  wire [2:0] _T_719 = _T_77 ? 3'h7 : _T_718;
  wire [2:0] _T_720 = _T_75 ? 3'h7 : _T_719;
  wire [2:0] _T_721 = _T_73 ? 3'h7 : _T_720;
  wire [2:0] _T_722 = _T_71 ? 3'h7 : _T_721;
  wire [2:0] _T_723 = _T_69 ? 3'h7 : _T_722;
  wire [2:0] _T_724 = _T_67 ? 3'h7 : _T_723;
  wire [2:0] _T_725 = _T_65 ? 3'h7 : _T_724;
  wire [2:0] _T_726 = _T_63 ? 3'h7 : _T_725;
  wire [2:0] _T_727 = _T_61 ? 3'h7 : _T_726;
  wire [2:0] _T_728 = _T_59 ? 3'h7 : _T_727;
  wire [2:0] _T_729 = _T_57 ? 3'h7 : _T_728;
  wire [2:0] _T_730 = _T_55 ? 3'h7 : _T_729;
  wire [2:0] _T_731 = _T_53 ? 3'h7 : _T_730;
  wire [2:0] _T_732 = _T_51 ? 3'h7 : _T_731;
  wire [2:0] _T_733 = _T_49 ? 3'h7 : _T_732;
  wire [2:0] _T_734 = _T_47 ? 3'h7 : _T_733;
  wire [2:0] _T_735 = _T_45 ? 3'h7 : _T_734;
  wire [2:0] _T_736 = _T_43 ? 3'h7 : _T_735;
  wire [2:0] _T_737 = _T_41 ? 3'h7 : _T_736;
  wire [2:0] _T_738 = _T_39 ? 3'h7 : _T_737;
  wire [2:0] _T_739 = _T_37 ? 3'h7 : _T_738;
  wire [2:0] c0_3 = _T_35 ? 3'h7 : _T_739;
  wire  _T_1220 = _T_99 ? 1'h0 : _T_101;
  wire  _T_1221 = _T_97 ? 1'h0 : _T_1220;
  wire  _T_1222 = _T_95 ? 1'h0 : _T_1221;
  wire  _T_1223 = _T_93 ? 1'h0 : _T_1222;
  wire  _T_1224 = _T_91 ? 1'h0 : _T_1223;
  wire  _T_1225 = _T_89 ? 1'h0 : _T_1224;
  wire  _T_1226 = _T_87 ? 1'h0 : _T_1225;
  wire  _T_1227 = _T_85 ? 1'h0 : _T_1226;
  wire  _T_1228 = _T_83 ? 1'h0 : _T_1227;
  wire  _T_1229 = _T_81 ? 1'h0 : _T_1228;
  wire  _T_1230 = _T_79 ? 1'h0 : _T_1229;
  wire  _T_1231 = _T_77 ? 1'h0 : _T_1230;
  wire  _T_1232 = _T_75 ? 1'h0 : _T_1231;
  wire  _T_1233 = _T_73 ? 1'h0 : _T_1232;
  wire  _T_1234 = _T_71 ? 1'h0 : _T_1233;
  wire  _T_1235 = _T_69 ? 1'h0 : _T_1234;
  wire  _T_1236 = _T_67 ? 1'h0 : _T_1235;
  wire  _T_1237 = _T_65 ? 1'h0 : _T_1236;
  wire  _T_1238 = _T_63 ? 1'h0 : _T_1237;
  wire  _T_1239 = _T_61 ? 1'h0 : _T_1238;
  wire  _T_1240 = _T_59 ? 1'h0 : _T_1239;
  wire  _T_1241 = _T_57 ? 1'h0 : _T_1240;
  wire  _T_1242 = _T_55 ? 1'h0 : _T_1241;
  wire  _T_1243 = _T_53 ? 1'h0 : _T_1242;
  wire  _T_1244 = _T_51 ? 1'h0 : _T_1243;
  wire  _T_1245 = _T_49 ? 1'h0 : _T_1244;
  wire  _T_1246 = _T_47 ? 1'h0 : _T_1245;
  wire  _T_1247 = _T_45 ? 1'h0 : _T_1246;
  wire  _T_1248 = _T_43 ? 1'h0 : _T_1247;
  wire  _T_1249 = _T_41 ? 1'h0 : _T_1248;
  wire  _T_1250 = _T_39 ? 1'h0 : _T_1249;
  wire  _T_1251 = _T_37 ? 1'h0 : _T_1250;
  wire  c0_11 = _T_35 ? 1'h0 : _T_1251;
  wire [4:0] _T_420 = _T_163 ? 5'h0 : 5'h13;
  wire [4:0] _T_421 = _T_161 ? 5'h0 : _T_420;
  wire [4:0] _T_422 = _T_159 ? 5'h0 : _T_421;
  wire [4:0] _T_423 = _T_157 ? 5'h0 : _T_422;
  wire [4:0] _T_424 = _T_155 ? 5'h0 : _T_423;
  wire [4:0] _T_425 = _T_153 ? 5'h0 : _T_424;
  wire [4:0] _T_426 = _T_151 ? 5'h0 : _T_425;
  wire [4:0] _T_427 = _T_149 ? 5'h0 : _T_426;
  wire [4:0] _T_428 = _T_147 ? 5'h0 : _T_427;
  wire [4:0] _T_429 = _T_145 ? 5'h13 : _T_428;
  wire [4:0] _T_430 = _T_143 ? 5'h13 : _T_429;
  wire [4:0] _T_431 = _T_141 ? 5'h0 : _T_430;
  wire [4:0] _T_432 = _T_139 ? 5'h0 : _T_431;
  wire [4:0] _T_433 = _T_137 ? 5'h0 : _T_432;
  wire [4:0] _T_434 = _T_135 ? 5'h0 : _T_433;
  wire [4:0] _T_435 = _T_133 ? 5'h0 : _T_434;
  wire [4:0] _T_436 = _T_131 ? 5'h0 : _T_435;
  wire [4:0] _T_437 = _T_129 ? 5'h0 : _T_436;
  wire [4:0] _T_438 = _T_127 ? 5'h0 : _T_437;
  wire [4:0] _T_439 = _T_125 ? 5'h0 : _T_438;
  wire [4:0] _T_440 = _T_123 ? 5'h0 : _T_439;
  wire [4:0] _T_441 = _T_121 ? 5'h0 : _T_440;
  wire [4:0] _T_442 = _T_119 ? 5'h0 : _T_441;
  wire [4:0] _T_443 = _T_117 ? 5'hb : _T_442;
  wire [4:0] _T_444 = _T_115 ? 5'h13 : _T_443;
  wire [4:0] _T_445 = _T_113 ? 5'h13 : _T_444;
  wire [4:0] _T_446 = _T_111 ? 5'h13 : _T_445;
  wire [4:0] _T_447 = _T_109 ? 5'h13 : _T_446;
  wire [4:0] _T_448 = _T_107 ? 5'h13 : _T_447;
  wire [4:0] _T_449 = _T_105 ? 5'h13 : _T_448;
  wire [4:0] _T_450 = _T_103 ? 5'h13 : _T_449;
  wire [4:0] _T_451 = _T_101 ? 5'h0 : _T_450;
  wire [4:0] _T_452 = _T_99 ? 5'h13 : _T_451;
  wire [4:0] _T_453 = _T_97 ? 5'h8 : _T_452;
  wire [4:0] _T_454 = _T_95 ? 5'h6 : _T_453;
  wire [4:0] _T_455 = _T_93 ? 5'h5 : _T_454;
  wire [4:0] _T_456 = _T_91 ? 5'h0 : _T_455;
  wire [4:0] _T_457 = _T_89 ? 5'ha : _T_456;
  wire [4:0] _T_458 = _T_87 ? 5'h9 : _T_457;
  wire [4:0] _T_459 = _T_85 ? 5'h4 : _T_458;
  wire [4:0] _T_460 = _T_83 ? 5'h3 : _T_459;
  wire [4:0] _T_461 = _T_81 ? 5'h2 : _T_460;
  wire [4:0] _T_462 = _T_79 ? 5'h13 : _T_461;
  wire [4:0] _T_463 = _T_77 ? 5'h13 : _T_462;
  wire [4:0] _T_464 = _T_75 ? 5'h11 : _T_463;
  wire [4:0] _T_465 = _T_73 ? 5'h12 : _T_464;
  wire [4:0] _T_466 = _T_71 ? 5'hf : _T_465;
  wire [4:0] _T_467 = _T_69 ? 5'h10 : _T_466;
  wire [4:0] _T_468 = _T_67 ? 5'he : _T_467;
  wire [4:0] _T_469 = _T_65 ? 5'hd : _T_468;
  wire [4:0] _T_470 = _T_63 ? 5'hc : _T_469;
  wire [4:0] _T_471 = _T_61 ? 5'h4 : _T_470;
  wire [4:0] _T_472 = _T_59 ? 5'h3 : _T_471;
  wire [4:0] _T_473 = _T_57 ? 5'h2 : _T_472;
  wire [4:0] _T_474 = _T_55 ? 5'h8 : _T_473;
  wire [4:0] _T_475 = _T_53 ? 5'h6 : _T_474;
  wire [4:0] _T_476 = _T_51 ? 5'h5 : _T_475;
  wire [4:0] _T_477 = _T_49 ? 5'h7 : _T_476;
  wire [4:0] _T_478 = _T_47 ? 5'ha : _T_477;
  wire [4:0] _T_479 = _T_45 ? 5'h9 : _T_478;
  wire [4:0] _T_480 = _T_43 ? 5'h1 : _T_479;
  wire [4:0] _T_481 = _T_41 ? 5'h0 : _T_480;
  wire [4:0] _T_482 = _T_39 ? 5'h13 : _T_481;
  wire [4:0] _T_483 = _T_37 ? 5'h13 : _T_482;
  wire [4:0] func = _T_35 ? 5'h13 : _T_483;
  wire  _aluOut_T = func == 5'h0;
  wire  _T_300 = _T_147 ? 1'h0 : _T_149 | (_T_151 | (_T_153 | (_T_155 | (_T_157 | (_T_159 | (_T_161 | _T_163))))));
  wire  _T_301 = _T_145 ? 1'h0 : _T_300;
  wire  _T_302 = _T_143 ? 1'h0 : _T_301;
  wire  _T_303 = _T_141 ? 1'h0 : _T_302;
  wire  _T_304 = _T_139 ? 1'h0 : _T_303;
  wire  _T_305 = _T_137 ? 1'h0 : _T_304;
  wire  _T_306 = _T_135 ? 1'h0 : _T_305;
  wire  _T_307 = _T_133 ? 1'h0 : _T_306;
  wire  _T_308 = _T_131 ? 1'h0 : _T_307;
  wire  _T_309 = _T_129 ? 1'h0 : _T_308;
  wire  _T_310 = _T_127 ? 1'h0 : _T_309;
  wire  _T_311 = _T_125 ? 1'h0 : _T_310;
  wire  _T_312 = _T_123 ? 1'h0 : _T_311;
  wire  _T_313 = _T_121 ? 1'h0 : _T_312;
  wire  _T_315 = _T_117 ? 1'h0 : _T_119 | _T_313;
  wire  _T_316 = _T_115 ? 1'h0 : _T_315;
  wire  _T_317 = _T_113 ? 1'h0 : _T_316;
  wire  _T_318 = _T_111 ? 1'h0 : _T_317;
  wire  _T_319 = _T_109 ? 1'h0 : _T_318;
  wire  _T_320 = _T_107 ? 1'h0 : _T_319;
  wire  _T_321 = _T_105 ? 1'h0 : _T_320;
  wire  _T_322 = _T_103 ? 1'h0 : _T_321;
  wire  _T_323 = _T_101 ? 1'h0 : _T_322;
  wire  _T_324 = _T_99 ? 1'h0 : _T_323;
  wire  _T_325 = _T_97 ? 1'h0 : _T_324;
  wire  _T_326 = _T_95 ? 1'h0 : _T_325;
  wire  _T_327 = _T_93 ? 1'h0 : _T_326;
  wire  _T_328 = _T_91 ? 1'h0 : _T_327;
  wire  _T_329 = _T_89 ? 1'h0 : _T_328;
  wire  _T_330 = _T_87 ? 1'h0 : _T_329;
  wire  _T_331 = _T_85 ? 1'h0 : _T_330;
  wire  _T_332 = _T_83 ? 1'h0 : _T_331;
  wire  _T_333 = _T_81 ? 1'h0 : _T_332;
  wire  _T_334 = _T_79 ? 1'h0 : _T_333;
  wire  _T_335 = _T_77 ? 1'h0 : _T_334;
  wire  _T_336 = _T_75 ? 1'h0 : _T_335;
  wire  _T_337 = _T_73 ? 1'h0 : _T_336;
  wire  _T_338 = _T_71 ? 1'h0 : _T_337;
  wire  _T_339 = _T_69 ? 1'h0 : _T_338;
  wire  _T_340 = _T_67 ? 1'h0 : _T_339;
  wire  _T_341 = _T_65 ? 1'h0 : _T_340;
  wire  _T_342 = _T_63 ? 1'h0 : _T_341;
  wire  _T_343 = _T_61 ? 1'h0 : _T_342;
  wire  _T_344 = _T_59 ? 1'h0 : _T_343;
  wire  _T_345 = _T_57 ? 1'h0 : _T_344;
  wire  _T_346 = _T_55 ? 1'h0 : _T_345;
  wire  _T_347 = _T_53 ? 1'h0 : _T_346;
  wire  _T_348 = _T_51 ? 1'h0 : _T_347;
  wire  _T_349 = _T_49 ? 1'h0 : _T_348;
  wire  _T_350 = _T_47 ? 1'h0 : _T_349;
  wire  _T_351 = _T_45 ? 1'h0 : _T_350;
  wire  _T_352 = _T_43 ? 1'h0 : _T_351;
  wire  _T_353 = _T_41 ? 1'h0 : _T_352;
  wire  _T_354 = _T_39 ? 1'h0 : _T_353;
  wire  _T_355 = _T_37 ? 1'h0 : _T_354;
  wire  op1Sel = _T_35 ? 1'h0 : _T_355;
  wire [4:0] j = inst[9:5];
  wire [31:0] rj = j == 5'h0 ? 32'h0 : GR_rj_MPORT_data;
  wire [31:0] aluOp1 = ~op1Sel ? rj : PC;
  wire [2:0] _T_356 = _T_163 ? 3'h5 : 3'h0;
  wire [2:0] _T_357 = _T_161 ? 3'h5 : _T_356;
  wire [2:0] _T_358 = _T_159 ? 3'h5 : _T_357;
  wire [2:0] _T_359 = _T_157 ? 3'h5 : _T_358;
  wire [2:0] _T_360 = _T_155 ? 3'h5 : _T_359;
  wire [2:0] _T_361 = _T_153 ? 3'h5 : _T_360;
  wire [2:0] _T_362 = _T_151 ? 3'h7 : _T_361;
  wire [2:0] _T_363 = _T_149 ? 3'h7 : _T_362;
  wire [2:0] _T_364 = _T_147 ? 3'h5 : _T_363;
  wire [2:0] _T_365 = _T_145 ? 3'h0 : _T_364;
  wire [2:0] _T_366 = _T_143 ? 3'h0 : _T_365;
  wire [2:0] _T_367 = _T_141 ? 3'h3 : _T_366;
  wire [2:0] _T_368 = _T_139 ? 3'h3 : _T_367;
  wire [2:0] _T_369 = _T_137 ? 3'h3 : _T_368;
  wire [2:0] _T_370 = _T_135 ? 3'h3 : _T_369;
  wire [2:0] _T_371 = _T_133 ? 3'h3 : _T_370;
  wire [2:0] _T_372 = _T_131 ? 3'h3 : _T_371;
  wire [2:0] _T_373 = _T_129 ? 3'h3 : _T_372;
  wire [2:0] _T_374 = _T_127 ? 3'h3 : _T_373;
  wire [2:0] _T_375 = _T_125 ? 3'h3 : _T_374;
  wire [2:0] _T_376 = _T_123 ? 3'h4 : _T_375;
  wire [2:0] _T_377 = _T_121 ? 3'h4 : _T_376;
  wire [2:0] _T_378 = _T_119 ? 3'h6 : _T_377;
  wire [2:0] _T_379 = _T_117 ? 3'h6 : _T_378;
  wire [2:0] _T_380 = _T_115 ? 3'h0 : _T_379;
  wire [2:0] _T_381 = _T_113 ? 3'h0 : _T_380;
  wire [2:0] _T_382 = _T_111 ? 3'h0 : _T_381;
  wire [2:0] _T_383 = _T_109 ? 3'h0 : _T_382;
  wire [2:0] _T_384 = _T_107 ? 3'h0 : _T_383;
  wire [2:0] _T_385 = _T_105 ? 3'h0 : _T_384;
  wire [2:0] _T_386 = _T_103 ? 3'h0 : _T_385;
  wire [2:0] _T_387 = _T_101 ? 3'h3 : _T_386;
  wire [2:0] _T_388 = _T_99 ? 3'h0 : _T_387;
  wire [2:0] _T_389 = _T_97 ? 3'h2 : _T_388;
  wire [2:0] _T_390 = _T_95 ? 3'h2 : _T_389;
  wire [2:0] _T_391 = _T_93 ? 3'h2 : _T_390;
  wire [2:0] _T_392 = _T_91 ? 3'h3 : _T_391;
  wire [2:0] _T_393 = _T_89 ? 3'h3 : _T_392;
  wire [2:0] _T_394 = _T_87 ? 3'h3 : _T_393;
  wire [2:0] _T_395 = _T_85 ? 3'h1 : _T_394;
  wire [2:0] _T_396 = _T_83 ? 3'h1 : _T_395;
  wire [2:0] _T_397 = _T_81 ? 3'h1 : _T_396;
  wire [2:0] _T_398 = _T_79 ? 3'h0 : _T_397;
  wire [2:0] _T_399 = _T_77 ? 3'h0 : _T_398;
  wire [2:0] _T_400 = _T_75 ? 3'h0 : _T_399;
  wire [2:0] _T_401 = _T_73 ? 3'h0 : _T_400;
  wire [2:0] _T_402 = _T_71 ? 3'h0 : _T_401;
  wire [2:0] _T_403 = _T_69 ? 3'h0 : _T_402;
  wire [2:0] _T_404 = _T_67 ? 3'h0 : _T_403;
  wire [2:0] _T_405 = _T_65 ? 3'h0 : _T_404;
  wire [2:0] _T_406 = _T_63 ? 3'h0 : _T_405;
  wire [2:0] _T_407 = _T_61 ? 3'h0 : _T_406;
  wire [2:0] _T_408 = _T_59 ? 3'h0 : _T_407;
  wire [2:0] _T_409 = _T_57 ? 3'h0 : _T_408;
  wire [2:0] _T_410 = _T_55 ? 3'h0 : _T_409;
  wire [2:0] _T_411 = _T_53 ? 3'h0 : _T_410;
  wire [2:0] _T_412 = _T_51 ? 3'h0 : _T_411;
  wire [2:0] _T_413 = _T_49 ? 3'h0 : _T_412;
  wire [2:0] _T_414 = _T_47 ? 3'h0 : _T_413;
  wire [2:0] _T_415 = _T_45 ? 3'h0 : _T_414;
  wire [2:0] _T_416 = _T_43 ? 3'h0 : _T_415;
  wire [2:0] _T_417 = _T_41 ? 3'h0 : _T_416;
  wire [2:0] _T_418 = _T_39 ? 3'h0 : _T_417;
  wire [2:0] _T_419 = _T_37 ? 3'h0 : _T_418;
  wire [2:0] op2Sel = _T_35 ? 3'h0 : _T_419;
  wire [3:0] _OFF26_T_2 = inst[9] ? 4'hf : 4'h0;
  wire [31:0] OFF26 = {_OFF26_T_2,inst[9:0],inst[25:10],2'h0};
  wire [31:0] UI20 = {inst[24:5],12'h0};
  wire [13:0] _OFF16_T_2 = inst[25] ? 14'h3fff : 14'h0;
  wire [31:0] OFF16 = {_OFF16_T_2,inst[25:10],2'h0};
  wire [17:0] _SI14_T_2 = inst[23] ? 18'h3ffff : 18'h0;
  wire [31:0] SI14 = {_SI14_T_2,inst[23:10]};
  wire [19:0] _SI12_T_2 = inst[21] ? 20'hfffff : 20'h0;
  wire [31:0] SI12 = {_SI12_T_2,inst[21:10]};
  wire [31:0] _aluOp2_WIRE_2 = {{20'd0}, inst[21:10]};
  wire [4:0] k = inst[14:10];
  wire [31:0] _aluOp2_WIRE_1 = {{27'd0}, k};
  wire  _T_773 = _T_97 ? 1'h0 : _T_99;
  wire  _T_774 = _T_95 ? 1'h0 : _T_773;
  wire  _T_775 = _T_93 ? 1'h0 : _T_774;
  wire  _T_776 = _T_91 ? 1'h0 : _T_775;
  wire  _T_777 = _T_89 ? 1'h0 : _T_776;
  wire  _T_778 = _T_87 ? 1'h0 : _T_777;
  wire  _T_779 = _T_85 ? 1'h0 : _T_778;
  wire  _T_780 = _T_83 ? 1'h0 : _T_779;
  wire  _T_781 = _T_81 ? 1'h0 : _T_780;
  wire  _T_782 = _T_79 ? 1'h0 : _T_781;
  wire  _T_783 = _T_77 ? 1'h0 : _T_782;
  wire  _T_784 = _T_75 ? 1'h0 : _T_783;
  wire  _T_785 = _T_73 ? 1'h0 : _T_784;
  wire  _T_786 = _T_71 ? 1'h0 : _T_785;
  wire  _T_787 = _T_69 ? 1'h0 : _T_786;
  wire  _T_788 = _T_67 ? 1'h0 : _T_787;
  wire  _T_789 = _T_65 ? 1'h0 : _T_788;
  wire  _T_790 = _T_63 ? 1'h0 : _T_789;
  wire  _T_791 = _T_61 ? 1'h0 : _T_790;
  wire  _T_792 = _T_59 ? 1'h0 : _T_791;
  wire  _T_793 = _T_57 ? 1'h0 : _T_792;
  wire  _T_794 = _T_55 ? 1'h0 : _T_793;
  wire  _T_795 = _T_53 ? 1'h0 : _T_794;
  wire  _T_796 = _T_51 ? 1'h0 : _T_795;
  wire  _T_797 = _T_49 ? 1'h0 : _T_796;
  wire  _T_798 = _T_47 ? 1'h0 : _T_797;
  wire  _T_799 = _T_45 ? 1'h0 : _T_798;
  wire  _T_800 = _T_43 ? 1'h0 : _T_799;
  wire  _T_801 = _T_41 ? 1'h0 : _T_800;
  wire  _T_802 = _T_39 ? 1'h0 : _T_801;
  wire  _T_803 = _T_37 ? 1'h0 : _T_802;
  wire  c0_4 = _T_35 ? 1'h0 : _T_803;
  wire [2:0] _T_1124 = _T_163 ? 3'h4 : 3'h0;
  wire [2:0] _T_1125 = _T_161 ? 3'h6 : _T_1124;
  wire [2:0] _T_1126 = _T_159 ? 3'h3 : _T_1125;
  wire [2:0] _T_1127 = _T_157 ? 3'h5 : _T_1126;
  wire [2:0] _T_1128 = _T_155 ? 3'h1 : _T_1127;
  wire [2:0] _T_1129 = _T_153 ? 3'h2 : _T_1128;
  wire [2:0] _T_1130 = _T_151 ? 3'h7 : _T_1129;
  wire [2:0] _T_1131 = _T_149 ? 3'h7 : _T_1130;
  wire [2:0] _T_1132 = _T_147 ? 3'h7 : _T_1131;
  wire [2:0] _T_1133 = _T_145 ? 3'h0 : _T_1132;
  wire [2:0] _T_1134 = _T_143 ? 3'h0 : _T_1133;
  wire [2:0] _T_1135 = _T_141 ? 3'h0 : _T_1134;
  wire [2:0] _T_1136 = _T_139 ? 3'h0 : _T_1135;
  wire [2:0] _T_1137 = _T_137 ? 3'h0 : _T_1136;
  wire [2:0] _T_1138 = _T_135 ? 3'h0 : _T_1137;
  wire [2:0] _T_1139 = _T_133 ? 3'h0 : _T_1138;
  wire [2:0] _T_1140 = _T_131 ? 3'h0 : _T_1139;
  wire [2:0] _T_1141 = _T_129 ? 3'h0 : _T_1140;
  wire [2:0] _T_1142 = _T_127 ? 3'h0 : _T_1141;
  wire [2:0] _T_1143 = _T_125 ? 3'h0 : _T_1142;
  wire [2:0] _T_1144 = _T_123 ? 3'h0 : _T_1143;
  wire [2:0] _T_1145 = _T_121 ? 3'h0 : _T_1144;
  wire [2:0] _T_1146 = _T_119 ? 3'h0 : _T_1145;
  wire [2:0] _T_1147 = _T_117 ? 3'h0 : _T_1146;
  wire [2:0] _T_1148 = _T_115 ? 3'h0 : _T_1147;
  wire [2:0] _T_1149 = _T_113 ? 3'h0 : _T_1148;
  wire [2:0] _T_1150 = _T_111 ? 3'h0 : _T_1149;
  wire [2:0] _T_1151 = _T_109 ? 3'h0 : _T_1150;
  wire [2:0] _T_1152 = _T_107 ? 3'h0 : _T_1151;
  wire [2:0] _T_1153 = _T_105 ? 3'h0 : _T_1152;
  wire [2:0] _T_1154 = _T_103 ? 3'h0 : _T_1153;
  wire [2:0] _T_1155 = _T_101 ? 3'h0 : _T_1154;
  wire [2:0] _T_1156 = _T_99 ? 3'h0 : _T_1155;
  wire [2:0] _T_1157 = _T_97 ? 3'h0 : _T_1156;
  wire [2:0] _T_1158 = _T_95 ? 3'h0 : _T_1157;
  wire [2:0] _T_1159 = _T_93 ? 3'h0 : _T_1158;
  wire [2:0] _T_1160 = _T_91 ? 3'h0 : _T_1159;
  wire [2:0] _T_1161 = _T_89 ? 3'h0 : _T_1160;
  wire [2:0] _T_1162 = _T_87 ? 3'h0 : _T_1161;
  wire [2:0] _T_1163 = _T_85 ? 3'h0 : _T_1162;
  wire [2:0] _T_1164 = _T_83 ? 3'h0 : _T_1163;
  wire [2:0] _T_1165 = _T_81 ? 3'h0 : _T_1164;
  wire [2:0] _T_1166 = _T_79 ? 3'h0 : _T_1165;
  wire [2:0] _T_1167 = _T_77 ? 3'h0 : _T_1166;
  wire [2:0] _T_1168 = _T_75 ? 3'h0 : _T_1167;
  wire [2:0] _T_1169 = _T_73 ? 3'h0 : _T_1168;
  wire [2:0] _T_1170 = _T_71 ? 3'h0 : _T_1169;
  wire [2:0] _T_1171 = _T_69 ? 3'h0 : _T_1170;
  wire [2:0] _T_1172 = _T_67 ? 3'h0 : _T_1171;
  wire [2:0] _T_1173 = _T_65 ? 3'h0 : _T_1172;
  wire [2:0] _T_1174 = _T_63 ? 3'h0 : _T_1173;
  wire [2:0] _T_1175 = _T_61 ? 3'h0 : _T_1174;
  wire [2:0] _T_1176 = _T_59 ? 3'h0 : _T_1175;
  wire [2:0] _T_1177 = _T_57 ? 3'h0 : _T_1176;
  wire [2:0] _T_1178 = _T_55 ? 3'h0 : _T_1177;
  wire [2:0] _T_1179 = _T_53 ? 3'h0 : _T_1178;
  wire [2:0] _T_1180 = _T_51 ? 3'h0 : _T_1179;
  wire [2:0] _T_1181 = _T_49 ? 3'h0 : _T_1180;
  wire [2:0] _T_1182 = _T_47 ? 3'h0 : _T_1181;
  wire [2:0] _T_1183 = _T_45 ? 3'h0 : _T_1182;
  wire [2:0] _T_1184 = _T_43 ? 3'h0 : _T_1183;
  wire [2:0] _T_1185 = _T_41 ? 3'h0 : _T_1184;
  wire [2:0] _T_1186 = _T_39 ? 3'h0 : _T_1185;
  wire [2:0] _T_1187 = _T_37 ? 3'h0 : _T_1186;
  wire [2:0] brType = _T_35 ? 3'h0 : _T_1187;
  wire  _kd_T_5 = ~(&c0_3[2:1]) | c0_4 | |brType;
  wire [4:0] kd = ~(&c0_3[2:1]) | c0_4 | |brType ? d : k;
  wire [31:0] rkd = kd == 5'h0 ? 32'h0 : GR_rkd_MPORT_data;
  wire [31:0] _GEN_71 = 3'h1 == op2Sel ? _aluOp2_WIRE_1 : rkd;
  wire [31:0] _GEN_72 = 3'h2 == op2Sel ? _aluOp2_WIRE_2 : _GEN_71;
  wire [31:0] _GEN_73 = 3'h3 == op2Sel ? SI12 : _GEN_72;
  wire [31:0] _GEN_74 = 3'h4 == op2Sel ? SI14 : _GEN_73;
  wire [31:0] _GEN_75 = 3'h5 == op2Sel ? OFF16 : _GEN_74;
  wire [31:0] _GEN_76 = 3'h6 == op2Sel ? UI20 : _GEN_75;
  wire [31:0] _GEN_77 = 3'h7 == op2Sel ? OFF26 : _GEN_76;
  wire [31:0] _aluOut_T_2 = aluOp1 + _GEN_77;
  wire [31:0] _aluOut_T_65 = _aluOut_T ? _aluOut_T_2 : 32'h0;
  wire  _aluOut_T_4 = func == 5'h1;
  wire [31:0] _aluOut_T_6 = aluOp1 - _GEN_77;
  wire [31:0] _aluOut_T_66 = _aluOut_T_4 ? _aluOut_T_6 : 32'h0;
  wire [31:0] _aluOut_T_84 = _aluOut_T_65 | _aluOut_T_66;
  wire  _aluOut_T_8 = func == 5'h2;
  wire [62:0] _GEN_7 = {{31'd0}, aluOp1};
  wire [62:0] _aluOut_T_10 = _GEN_7 << _GEN_77[4:0];
  wire [31:0] _aluOut_T_67 = _aluOut_T_8 ? _aluOut_T_10[31:0] : 32'h0;
  wire [31:0] _aluOut_T_85 = _aluOut_T_84 | _aluOut_T_67;
  wire  _aluOut_T_12 = func == 5'h3;
  wire [31:0] _aluOut_T_14 = aluOp1 >> _GEN_77[4:0];
  wire [31:0] _aluOut_T_68 = _aluOut_T_12 ? _aluOut_T_14 : 32'h0;
  wire [31:0] _aluOut_T_86 = _aluOut_T_85 | _aluOut_T_68;
  wire  _aluOut_T_16 = func == 5'h4;
  wire [31:0] aluOut_sa = ~op1Sel ? rj : PC;
  wire [31:0] _aluOut_T_19 = $signed(aluOut_sa) >>> _GEN_77[4:0];
  wire [31:0] _aluOut_T_69 = _aluOut_T_16 ? _aluOut_T_19 : 32'h0;
  wire [31:0] _aluOut_T_87 = _aluOut_T_86 | _aluOut_T_69;
  wire  _aluOut_T_21 = func == 5'h5;
  wire [31:0] _aluOut_T_22 = aluOp1 & _GEN_77;
  wire [31:0] _aluOut_T_70 = _aluOut_T_21 ? _aluOut_T_22 : 32'h0;
  wire [31:0] _aluOut_T_88 = _aluOut_T_87 | _aluOut_T_70;
  wire  _aluOut_T_24 = func == 5'h6;
  wire [31:0] _aluOut_T_25 = aluOp1 | _GEN_77;
  wire [31:0] _aluOut_T_71 = _aluOut_T_24 ? _aluOut_T_25 : 32'h0;
  wire [31:0] _aluOut_T_89 = _aluOut_T_88 | _aluOut_T_71;
  wire  _aluOut_T_27 = func == 5'h7;
  wire [31:0] _aluOut_T_29 = ~_aluOut_T_25;
  wire [31:0] _aluOut_T_72 = _aluOut_T_27 ? _aluOut_T_29 : 32'h0;
  wire [31:0] _aluOut_T_90 = _aluOut_T_89 | _aluOut_T_72;
  wire  _aluOut_T_31 = func == 5'h8;
  wire [31:0] _aluOut_T_32 = aluOp1 ^ _GEN_77;
  wire [31:0] _aluOut_T_73 = _aluOut_T_31 ? _aluOut_T_32 : 32'h0;
  wire [31:0] _aluOut_T_91 = _aluOut_T_90 | _aluOut_T_73;
  wire  _aluOut_T_34 = func == 5'h9;
  wire [31:0] aluOut_sb = 3'h7 == op2Sel ? OFF26 : _GEN_76;
  wire  _aluOut_T_35 = $signed(aluOut_sa) < $signed(aluOut_sb);
  wire  _aluOut_T_74 = _aluOut_T_34 & _aluOut_T_35;
  wire [31:0] _GEN_2357 = {{31'd0}, _aluOut_T_74};
  wire [31:0] _aluOut_T_92 = _aluOut_T_91 | _GEN_2357;
  wire  _aluOut_T_36 = func == 5'ha;
  wire  _aluOut_T_37 = aluOp1 < _GEN_77;
  wire  _aluOut_T_75 = _aluOut_T_36 & _aluOut_T_37;
  wire [31:0] _GEN_2358 = {{31'd0}, _aluOut_T_75};
  wire [31:0] _aluOut_T_93 = _aluOut_T_92 | _GEN_2358;
  wire  _aluOut_T_38 = func == 5'hb;
  wire [31:0] _aluOut_T_76 = _aluOut_T_38 ? _GEN_77 : 32'h0;
  wire [31:0] _aluOut_T_94 = _aluOut_T_93 | _aluOut_T_76;
  wire  _aluOut_T_40 = func == 5'hc;
  wire [63:0] _aluOut_T_42 = $signed(aluOut_sa) * $signed(aluOut_sb);
  wire [31:0] _aluOut_T_77 = _aluOut_T_40 ? _aluOut_T_42[31:0] : 32'h0;
  wire [31:0] _aluOut_T_95 = _aluOut_T_94 | _aluOut_T_77;
  wire  _aluOut_T_44 = func == 5'hd;
  wire [31:0] _aluOut_T_78 = _aluOut_T_44 ? _aluOut_T_42[63:32] : 32'h0;
  wire [31:0] _aluOut_T_96 = _aluOut_T_95 | _aluOut_T_78;
  wire  _aluOut_T_48 = func == 5'he;
  wire [63:0] _aluOut_T_49 = aluOp1 * _GEN_77;
  wire [31:0] _aluOut_T_79 = _aluOut_T_48 ? _aluOut_T_49[63:32] : 32'h0;
  wire [31:0] _aluOut_T_97 = _aluOut_T_96 | _aluOut_T_79;
  wire  _aluOut_T_51 = func == 5'hf;
  wire [31:0] _aluOut_T_53 = $signed(aluOut_sa) % $signed(aluOut_sb);
  wire [31:0] _aluOut_T_80 = _aluOut_T_51 ? _aluOut_T_53 : 32'h0;
  wire [31:0] _aluOut_T_98 = _aluOut_T_97 | _aluOut_T_80;
  wire  _aluOut_T_55 = func == 5'h10;
  wire [32:0] _aluOut_T_57 = $signed(aluOut_sa) / $signed(aluOut_sb);
  wire [31:0] _aluOut_T_81 = _aluOut_T_55 ? _aluOut_T_57[31:0] : 32'h0;
  wire [31:0] _aluOut_T_99 = _aluOut_T_98 | _aluOut_T_81;
  wire  _aluOut_T_59 = func == 5'h11;
  wire [31:0] _aluOut_T_60 = aluOp1 % _GEN_77;
  wire [31:0] _aluOut_T_82 = _aluOut_T_59 ? _aluOut_T_60 : 32'h0;
  wire [31:0] _aluOut_T_100 = _aluOut_T_99 | _aluOut_T_82;
  wire  _aluOut_T_62 = func == 5'h12;
  wire [31:0] _aluOut_T_63 = aluOp1 / _GEN_77;
  wire [31:0] _aluOut_T_83 = _aluOut_T_62 ? _aluOut_T_63 : 32'h0;
  wire [31:0] aluOut = _aluOut_T_100 | _aluOut_T_83;
  wire  memALE = aluOut[0] & c0_3[2:1] == 2'h1 | |aluOut[1:0] & c0_3[2:1] == 2'h2;
  wire  _EXVA_T = c0_3 != 3'h7;
  wire [31:0] _EXVA_T_4 = _EXVA_T ? aluOut : 32'h0;
  wire  _EXVA_T_1 = c0_7 == 3'h1;
  wire [31:0] _EXVA_T_2 = {csrs_9_VPPN,13'h0};
  wire [31:0] _EXVA_T_5 = _EXVA_T_1 ? _EXVA_T_2 : 32'h0;
  wire [31:0] _EXVA_T_7 = _EXVA_T_4 | _EXVA_T_5;
  wire [31:0] _EXVA_T_6 = _INE_T_1 ? rkd : 32'h0;
  wire [31:0] EXVA = _EXVA_T_7 | _EXVA_T_6;
  wire  vaMatch_0_1 = tlb_0_VPPN[18:9] == EXVA[31:22] & (tlb_0_PS == 6'h15 | tlb_0_VPPN[8:0] == EXVA[21:13]);
  wire [9:0] EXASID = _INE_T_1 ? rj[9:0] : asid_ASID;
  wire  asidMatch_0_1 = tlb_0_ASID == EXASID;
  wire  tlbHit_0_1 = tlb_0_E & vaMatch_0_1 & (tlb_0_G | asidMatch_0_1);
  wire  vaMatch_1_1 = tlb_1_VPPN[18:9] == EXVA[31:22] & (tlb_1_PS == 6'h15 | tlb_1_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_1_1 = tlb_1_ASID == EXASID;
  wire  tlbHit_1_1 = tlb_1_E & vaMatch_1_1 & (tlb_1_G | asidMatch_1_1);
  wire  vaMatch_2_1 = tlb_2_VPPN[18:9] == EXVA[31:22] & (tlb_2_PS == 6'h15 | tlb_2_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_2_1 = tlb_2_ASID == EXASID;
  wire  tlbHit_2_1 = tlb_2_E & vaMatch_2_1 & (tlb_2_G | asidMatch_2_1);
  wire  vaMatch_3_1 = tlb_3_VPPN[18:9] == EXVA[31:22] & (tlb_3_PS == 6'h15 | tlb_3_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_3_1 = tlb_3_ASID == EXASID;
  wire  tlbHit_3_1 = tlb_3_E & vaMatch_3_1 & (tlb_3_G | asidMatch_3_1);
  wire  vaMatch_4_1 = tlb_4_VPPN[18:9] == EXVA[31:22] & (tlb_4_PS == 6'h15 | tlb_4_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_4_1 = tlb_4_ASID == EXASID;
  wire  tlbHit_4_1 = tlb_4_E & vaMatch_4_1 & (tlb_4_G | asidMatch_4_1);
  wire  vaMatch_5_1 = tlb_5_VPPN[18:9] == EXVA[31:22] & (tlb_5_PS == 6'h15 | tlb_5_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_5_1 = tlb_5_ASID == EXASID;
  wire  tlbHit_5_1 = tlb_5_E & vaMatch_5_1 & (tlb_5_G | asidMatch_5_1);
  wire  vaMatch_6_1 = tlb_6_VPPN[18:9] == EXVA[31:22] & (tlb_6_PS == 6'h15 | tlb_6_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_6_1 = tlb_6_ASID == EXASID;
  wire  tlbHit_6_1 = tlb_6_E & vaMatch_6_1 & (tlb_6_G | asidMatch_6_1);
  wire  vaMatch_7_1 = tlb_7_VPPN[18:9] == EXVA[31:22] & (tlb_7_PS == 6'h15 | tlb_7_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_7_1 = tlb_7_ASID == EXASID;
  wire  tlbHit_7_1 = tlb_7_E & vaMatch_7_1 & (tlb_7_G | asidMatch_7_1);
  wire  vaMatch_8_1 = tlb_8_VPPN[18:9] == EXVA[31:22] & (tlb_8_PS == 6'h15 | tlb_8_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_8_1 = tlb_8_ASID == EXASID;
  wire  tlbHit_8_1 = tlb_8_E & vaMatch_8_1 & (tlb_8_G | asidMatch_8_1);
  wire  vaMatch_9_1 = tlb_9_VPPN[18:9] == EXVA[31:22] & (tlb_9_PS == 6'h15 | tlb_9_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_9_1 = tlb_9_ASID == EXASID;
  wire  tlbHit_9_1 = tlb_9_E & vaMatch_9_1 & (tlb_9_G | asidMatch_9_1);
  wire  vaMatch_10_1 = tlb_10_VPPN[18:9] == EXVA[31:22] & (tlb_10_PS == 6'h15 | tlb_10_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_10_1 = tlb_10_ASID == EXASID;
  wire  tlbHit_10_1 = tlb_10_E & vaMatch_10_1 & (tlb_10_G | asidMatch_10_1);
  wire  vaMatch_11_1 = tlb_11_VPPN[18:9] == EXVA[31:22] & (tlb_11_PS == 6'h15 | tlb_11_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_11_1 = tlb_11_ASID == EXASID;
  wire  tlbHit_11_1 = tlb_11_E & vaMatch_11_1 & (tlb_11_G | asidMatch_11_1);
  wire  vaMatch_12_1 = tlb_12_VPPN[18:9] == EXVA[31:22] & (tlb_12_PS == 6'h15 | tlb_12_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_12_1 = tlb_12_ASID == EXASID;
  wire  tlbHit_12_1 = tlb_12_E & vaMatch_12_1 & (tlb_12_G | asidMatch_12_1);
  wire  vaMatch_13_1 = tlb_13_VPPN[18:9] == EXVA[31:22] & (tlb_13_PS == 6'h15 | tlb_13_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_13_1 = tlb_13_ASID == EXASID;
  wire  tlbHit_13_1 = tlb_13_E & vaMatch_13_1 & (tlb_13_G | asidMatch_13_1);
  wire  vaMatch_14_1 = tlb_14_VPPN[18:9] == EXVA[31:22] & (tlb_14_PS == 6'h15 | tlb_14_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_14_1 = tlb_14_ASID == EXASID;
  wire  tlbHit_14_1 = tlb_14_E & vaMatch_14_1 & (tlb_14_G | asidMatch_14_1);
  wire  vaMatch_15_1 = tlb_15_VPPN[18:9] == EXVA[31:22] & (tlb_15_PS == 6'h15 | tlb_15_VPPN[8:0] == EXVA[21:13]);
  wire  asidMatch_15_1 = tlb_15_ASID == EXASID;
  wire  tlbHit_15_1 = tlb_15_E & vaMatch_15_1 & (tlb_15_G | asidMatch_15_1);
  wire  _miss_T_30 = tlbHit_0_1 | tlbHit_1_1 | tlbHit_2_1 | tlbHit_3_1 | tlbHit_4_1 | tlbHit_5_1 | tlbHit_6_1 |
    tlbHit_7_1 | tlbHit_8_1 | tlbHit_9_1 | tlbHit_10_1 | tlbHit_11_1 | tlbHit_12_1 | tlbHit_13_1 | tlbHit_14_1 |
    tlbHit_15_1;
  wire  _GEN_81 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : ~(tlbHit_0_1 |
    tlbHit_1_1 | tlbHit_2_1 | tlbHit_3_1 | tlbHit_4_1 | tlbHit_5_1 | tlbHit_6_1 | tlbHit_7_1 | tlbHit_8_1 | tlbHit_9_1
     | tlbHit_10_1 | tlbHit_11_1 | tlbHit_12_1 | tlbHit_13_1 | tlbHit_14_1 | tlbHit_15_1);
  wire  miss_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_81;
  wire  _T_1264 = _T_139 ? 1'h0 : _T_141;
  wire  _T_1265 = _T_137 ? 1'h0 : _T_1264;
  wire  _T_1266 = _T_135 ? 1'h0 : _T_1265;
  wire  _T_1267 = _T_133 ? 1'h0 : _T_1266;
  wire  _T_1268 = _T_131 ? 1'h0 : _T_1267;
  wire  _T_1269 = _T_129 ? 1'h0 : _T_1268;
  wire  _T_1270 = _T_127 ? 1'h0 : _T_1269;
  wire  _T_1271 = _T_125 ? 1'h0 : _T_1270;
  wire  _T_1272 = _T_123 ? 1'h0 : _T_1271;
  wire  _T_1273 = _T_121 ? 1'h0 : _T_1272;
  wire  _T_1274 = _T_119 ? 1'h0 : _T_1273;
  wire  _T_1275 = _T_117 ? 1'h0 : _T_1274;
  wire  _T_1276 = _T_115 ? 1'h0 : _T_1275;
  wire  _T_1277 = _T_113 ? 1'h0 : _T_1276;
  wire  _T_1278 = _T_111 ? 1'h0 : _T_1277;
  wire  _T_1279 = _T_109 ? 1'h0 : _T_1278;
  wire  _T_1280 = _T_107 ? 1'h0 : _T_1279;
  wire  _T_1281 = _T_105 ? 1'h0 : _T_1280;
  wire  _T_1282 = _T_103 ? 1'h0 : _T_1281;
  wire  _T_1283 = _T_101 ? 1'h0 : _T_1282;
  wire  _T_1284 = _T_99 ? 1'h0 : _T_1283;
  wire  _T_1285 = _T_97 ? 1'h0 : _T_1284;
  wire  _T_1286 = _T_95 ? 1'h0 : _T_1285;
  wire  _T_1287 = _T_93 ? 1'h0 : _T_1286;
  wire  _T_1288 = _T_91 ? 1'h0 : _T_1287;
  wire  _T_1289 = _T_89 ? 1'h0 : _T_1288;
  wire  _T_1290 = _T_87 ? 1'h0 : _T_1289;
  wire  _T_1291 = _T_85 ? 1'h0 : _T_1290;
  wire  _T_1292 = _T_83 ? 1'h0 : _T_1291;
  wire  _T_1293 = _T_81 ? 1'h0 : _T_1292;
  wire  _T_1294 = _T_79 ? 1'h0 : _T_1293;
  wire  _T_1295 = _T_77 ? 1'h0 : _T_1294;
  wire  _T_1296 = _T_75 ? 1'h0 : _T_1295;
  wire  _T_1297 = _T_73 ? 1'h0 : _T_1296;
  wire  _T_1298 = _T_71 ? 1'h0 : _T_1297;
  wire  _T_1299 = _T_69 ? 1'h0 : _T_1298;
  wire  _T_1300 = _T_67 ? 1'h0 : _T_1299;
  wire  _T_1301 = _T_65 ? 1'h0 : _T_1300;
  wire  _T_1302 = _T_63 ? 1'h0 : _T_1301;
  wire  _T_1303 = _T_61 ? 1'h0 : _T_1302;
  wire  _T_1304 = _T_59 ? 1'h0 : _T_1303;
  wire  _T_1305 = _T_57 ? 1'h0 : _T_1304;
  wire  _T_1306 = _T_55 ? 1'h0 : _T_1305;
  wire  _T_1307 = _T_53 ? 1'h0 : _T_1306;
  wire  _T_1308 = _T_51 ? 1'h0 : _T_1307;
  wire  _T_1309 = _T_49 ? 1'h0 : _T_1308;
  wire  _T_1310 = _T_47 ? 1'h0 : _T_1309;
  wire  _T_1311 = _T_45 ? 1'h0 : _T_1310;
  wire  _T_1312 = _T_43 ? 1'h0 : _T_1311;
  wire  _T_1313 = _T_41 ? 1'h0 : _T_1312;
  wire  _T_1314 = _T_39 ? 1'h0 : _T_1313;
  wire  _T_1315 = _T_37 ? 1'h0 : _T_1314;
  wire  c0_12 = _T_35 ? 1'h0 : _T_1315;
  wire  _TLBR_T = ~c0_12;
  wire  _GEN_112 = miss_1 ? ~c0_12 : _GEN_56;
  wire  _GEN_129 = crmd_DA ? _GEN_56 : _GEN_112;
  wire  _GEN_138 = memALE ? _GEN_56 : _GEN_129;
  wire  _GEN_147 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? _GEN_56 : _GEN_138;
  wire  _GEN_159 = ID_OK ? _GEN_147 : _GEN_56;
  wire  TLBR = dStallReg ? _GEN_56 : _GEN_159;
  wire  _GEN_135 = memALE & _TLBR_T;
  wire  _GEN_145 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_135;
  wire  _GEN_157 = ID_OK & _GEN_145;
  wire  ALE = dStallReg ? 1'h0 : _GEN_157;
  wire [7:0] excp_lo = {ALE,SYS,BRK,INE,2'h0,1'h0,TLBR};
  wire  _GEN_47 = ~INT & ~idle & _T_31;
  wire  ADEF = dStallReg | iStallReg ? 1'h0 : _GEN_47;
  wire [5:0] _foundTLB_T_868 = tlbHit_0_1 ? tlb_0_PS : 6'h0;
  wire [5:0] _foundTLB_T_869 = tlbHit_1_1 ? tlb_1_PS : 6'h0;
  wire [5:0] _foundTLB_T_884 = _foundTLB_T_868 | _foundTLB_T_869;
  wire [5:0] _foundTLB_T_870 = tlbHit_2_1 ? tlb_2_PS : 6'h0;
  wire [5:0] _foundTLB_T_885 = _foundTLB_T_884 | _foundTLB_T_870;
  wire [5:0] _foundTLB_T_871 = tlbHit_3_1 ? tlb_3_PS : 6'h0;
  wire [5:0] _foundTLB_T_886 = _foundTLB_T_885 | _foundTLB_T_871;
  wire [5:0] _foundTLB_T_872 = tlbHit_4_1 ? tlb_4_PS : 6'h0;
  wire [5:0] _foundTLB_T_887 = _foundTLB_T_886 | _foundTLB_T_872;
  wire [5:0] _foundTLB_T_873 = tlbHit_5_1 ? tlb_5_PS : 6'h0;
  wire [5:0] _foundTLB_T_888 = _foundTLB_T_887 | _foundTLB_T_873;
  wire [5:0] _foundTLB_T_874 = tlbHit_6_1 ? tlb_6_PS : 6'h0;
  wire [5:0] _foundTLB_T_889 = _foundTLB_T_888 | _foundTLB_T_874;
  wire [5:0] _foundTLB_T_875 = tlbHit_7_1 ? tlb_7_PS : 6'h0;
  wire [5:0] _foundTLB_T_890 = _foundTLB_T_889 | _foundTLB_T_875;
  wire [5:0] _foundTLB_T_876 = tlbHit_8_1 ? tlb_8_PS : 6'h0;
  wire [5:0] _foundTLB_T_891 = _foundTLB_T_890 | _foundTLB_T_876;
  wire [5:0] _foundTLB_T_877 = tlbHit_9_1 ? tlb_9_PS : 6'h0;
  wire [5:0] _foundTLB_T_892 = _foundTLB_T_891 | _foundTLB_T_877;
  wire [5:0] _foundTLB_T_878 = tlbHit_10_1 ? tlb_10_PS : 6'h0;
  wire [5:0] _foundTLB_T_893 = _foundTLB_T_892 | _foundTLB_T_878;
  wire [5:0] _foundTLB_T_879 = tlbHit_11_1 ? tlb_11_PS : 6'h0;
  wire [5:0] _foundTLB_T_894 = _foundTLB_T_893 | _foundTLB_T_879;
  wire [5:0] _foundTLB_T_880 = tlbHit_12_1 ? tlb_12_PS : 6'h0;
  wire [5:0] _foundTLB_T_895 = _foundTLB_T_894 | _foundTLB_T_880;
  wire [5:0] _foundTLB_T_881 = tlbHit_13_1 ? tlb_13_PS : 6'h0;
  wire [5:0] _foundTLB_T_896 = _foundTLB_T_895 | _foundTLB_T_881;
  wire [5:0] _foundTLB_T_882 = tlbHit_14_1 ? tlb_14_PS : 6'h0;
  wire [5:0] _foundTLB_T_897 = _foundTLB_T_896 | _foundTLB_T_882;
  wire [5:0] _foundTLB_T_883 = tlbHit_15_1 ? tlb_15_PS : 6'h0;
  wire [5:0] foundTLB_1_PS = _foundTLB_T_897 | _foundTLB_T_883;
  wire  _oddPG_T_3 = foundTLB_1_PS == 6'hc;
  wire  oddPG_1 = foundTLB_1_PS == 6'hc ? EXVA[12] : EXVA[21];
  wire  _foundTLB_T_480 = tlbHit_15_1 & tlb_15_P1_V;
  wire  foundTLB_1_P1_V = tlbHit_0_1 & tlb_0_P1_V | tlbHit_1_1 & tlb_1_P1_V | tlbHit_2_1 & tlb_2_P1_V | tlbHit_3_1 &
    tlb_3_P1_V | tlbHit_4_1 & tlb_4_P1_V | tlbHit_5_1 & tlb_5_P1_V | tlbHit_6_1 & tlb_6_P1_V | tlbHit_7_1 & tlb_7_P1_V
     | tlbHit_8_1 & tlb_8_P1_V | tlbHit_9_1 & tlb_9_P1_V | tlbHit_10_1 & tlb_10_P1_V | tlbHit_11_1 & tlb_11_P1_V |
    tlbHit_12_1 & tlb_12_P1_V | tlbHit_13_1 & tlb_13_P1_V | tlbHit_14_1 & tlb_14_P1_V | _foundTLB_T_480;
  wire  _foundTLB_T_635 = tlbHit_15_1 & tlb_15_P0_V;
  wire  foundTLB_1_P0_V = tlbHit_0_1 & tlb_0_P0_V | tlbHit_1_1 & tlb_1_P0_V | tlbHit_2_1 & tlb_2_P0_V | tlbHit_3_1 &
    tlb_3_P0_V | tlbHit_4_1 & tlb_4_P0_V | tlbHit_5_1 & tlb_5_P0_V | tlbHit_6_1 & tlb_6_P0_V | tlbHit_7_1 & tlb_7_P0_V
     | tlbHit_8_1 & tlb_8_P0_V | tlbHit_9_1 & tlb_9_P0_V | tlbHit_10_1 & tlb_10_P0_V | tlbHit_11_1 & tlb_11_P0_V |
    tlbHit_12_1 & tlb_12_P0_V | tlbHit_13_1 & tlb_13_P0_V | tlbHit_14_1 & tlb_14_P0_V | _foundTLB_T_635;
  wire  foundP_1_V = oddPG_1 ? foundTLB_1_P1_V : foundTLB_1_P0_V;
  wire  _GEN_82 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : ~foundP_1_V;
  wire  invalid_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_82;
  wire [1:0] _foundTLB_T_558 = tlbHit_0_1 ? tlb_0_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_559 = tlbHit_1_1 ? tlb_1_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_574 = _foundTLB_T_558 | _foundTLB_T_559;
  wire [1:0] _foundTLB_T_560 = tlbHit_2_1 ? tlb_2_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_575 = _foundTLB_T_574 | _foundTLB_T_560;
  wire [1:0] _foundTLB_T_561 = tlbHit_3_1 ? tlb_3_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_576 = _foundTLB_T_575 | _foundTLB_T_561;
  wire [1:0] _foundTLB_T_562 = tlbHit_4_1 ? tlb_4_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_577 = _foundTLB_T_576 | _foundTLB_T_562;
  wire [1:0] _foundTLB_T_563 = tlbHit_5_1 ? tlb_5_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_578 = _foundTLB_T_577 | _foundTLB_T_563;
  wire [1:0] _foundTLB_T_564 = tlbHit_6_1 ? tlb_6_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_579 = _foundTLB_T_578 | _foundTLB_T_564;
  wire [1:0] _foundTLB_T_565 = tlbHit_7_1 ? tlb_7_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_580 = _foundTLB_T_579 | _foundTLB_T_565;
  wire [1:0] _foundTLB_T_566 = tlbHit_8_1 ? tlb_8_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_581 = _foundTLB_T_580 | _foundTLB_T_566;
  wire [1:0] _foundTLB_T_567 = tlbHit_9_1 ? tlb_9_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_582 = _foundTLB_T_581 | _foundTLB_T_567;
  wire [1:0] _foundTLB_T_568 = tlbHit_10_1 ? tlb_10_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_583 = _foundTLB_T_582 | _foundTLB_T_568;
  wire [1:0] _foundTLB_T_569 = tlbHit_11_1 ? tlb_11_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_584 = _foundTLB_T_583 | _foundTLB_T_569;
  wire [1:0] _foundTLB_T_570 = tlbHit_12_1 ? tlb_12_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_585 = _foundTLB_T_584 | _foundTLB_T_570;
  wire [1:0] _foundTLB_T_571 = tlbHit_13_1 ? tlb_13_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_586 = _foundTLB_T_585 | _foundTLB_T_571;
  wire [1:0] _foundTLB_T_572 = tlbHit_14_1 ? tlb_14_P1_PLV : 2'h0;
  wire [1:0] _foundTLB_T_587 = _foundTLB_T_586 | _foundTLB_T_572;
  wire [1:0] _foundTLB_T_573 = tlbHit_15_1 ? tlb_15_P1_PLV : 2'h0;
  wire [1:0] foundTLB_1_P1_PLV = _foundTLB_T_587 | _foundTLB_T_573;
  wire [1:0] _foundTLB_T_713 = tlbHit_0_1 ? tlb_0_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_714 = tlbHit_1_1 ? tlb_1_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_729 = _foundTLB_T_713 | _foundTLB_T_714;
  wire [1:0] _foundTLB_T_715 = tlbHit_2_1 ? tlb_2_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_730 = _foundTLB_T_729 | _foundTLB_T_715;
  wire [1:0] _foundTLB_T_716 = tlbHit_3_1 ? tlb_3_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_731 = _foundTLB_T_730 | _foundTLB_T_716;
  wire [1:0] _foundTLB_T_717 = tlbHit_4_1 ? tlb_4_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_732 = _foundTLB_T_731 | _foundTLB_T_717;
  wire [1:0] _foundTLB_T_718 = tlbHit_5_1 ? tlb_5_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_733 = _foundTLB_T_732 | _foundTLB_T_718;
  wire [1:0] _foundTLB_T_719 = tlbHit_6_1 ? tlb_6_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_734 = _foundTLB_T_733 | _foundTLB_T_719;
  wire [1:0] _foundTLB_T_720 = tlbHit_7_1 ? tlb_7_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_735 = _foundTLB_T_734 | _foundTLB_T_720;
  wire [1:0] _foundTLB_T_721 = tlbHit_8_1 ? tlb_8_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_736 = _foundTLB_T_735 | _foundTLB_T_721;
  wire [1:0] _foundTLB_T_722 = tlbHit_9_1 ? tlb_9_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_737 = _foundTLB_T_736 | _foundTLB_T_722;
  wire [1:0] _foundTLB_T_723 = tlbHit_10_1 ? tlb_10_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_738 = _foundTLB_T_737 | _foundTLB_T_723;
  wire [1:0] _foundTLB_T_724 = tlbHit_11_1 ? tlb_11_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_739 = _foundTLB_T_738 | _foundTLB_T_724;
  wire [1:0] _foundTLB_T_725 = tlbHit_12_1 ? tlb_12_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_740 = _foundTLB_T_739 | _foundTLB_T_725;
  wire [1:0] _foundTLB_T_726 = tlbHit_13_1 ? tlb_13_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_741 = _foundTLB_T_740 | _foundTLB_T_726;
  wire [1:0] _foundTLB_T_727 = tlbHit_14_1 ? tlb_14_P0_PLV : 2'h0;
  wire [1:0] _foundTLB_T_742 = _foundTLB_T_741 | _foundTLB_T_727;
  wire [1:0] _foundTLB_T_728 = tlbHit_15_1 ? tlb_15_P0_PLV : 2'h0;
  wire [1:0] foundTLB_1_P0_PLV = _foundTLB_T_742 | _foundTLB_T_728;
  wire [1:0] foundP_1_PLV = oddPG_1 ? foundTLB_1_P1_PLV : foundTLB_1_P0_PLV;
  wire  _GEN_83 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : crmd_PLV >
    foundP_1_PLV;
  wire  ppi_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_83;
  reg  tlb_0_P1_D;
  reg  tlb_1_P1_D;
  reg  tlb_2_P1_D;
  reg  tlb_3_P1_D;
  reg  tlb_4_P1_D;
  reg  tlb_5_P1_D;
  reg  tlb_6_P1_D;
  reg  tlb_7_P1_D;
  reg  tlb_8_P1_D;
  reg  tlb_9_P1_D;
  reg  tlb_10_P1_D;
  reg  tlb_11_P1_D;
  reg  tlb_12_P1_D;
  reg  tlb_13_P1_D;
  reg  tlb_14_P1_D;
  reg  tlb_15_P1_D;
  wire  _foundTLB_T_511 = tlbHit_15_1 & tlb_15_P1_D;
  wire  foundTLB_1_P1_D = tlbHit_0_1 & tlb_0_P1_D | tlbHit_1_1 & tlb_1_P1_D | tlbHit_2_1 & tlb_2_P1_D | tlbHit_3_1 &
    tlb_3_P1_D | tlbHit_4_1 & tlb_4_P1_D | tlbHit_5_1 & tlb_5_P1_D | tlbHit_6_1 & tlb_6_P1_D | tlbHit_7_1 & tlb_7_P1_D
     | tlbHit_8_1 & tlb_8_P1_D | tlbHit_9_1 & tlb_9_P1_D | tlbHit_10_1 & tlb_10_P1_D | tlbHit_11_1 & tlb_11_P1_D |
    tlbHit_12_1 & tlb_12_P1_D | tlbHit_13_1 & tlb_13_P1_D | tlbHit_14_1 & tlb_14_P1_D | _foundTLB_T_511;
  reg  tlb_0_P0_D;
  reg  tlb_1_P0_D;
  reg  tlb_2_P0_D;
  reg  tlb_3_P0_D;
  reg  tlb_4_P0_D;
  reg  tlb_5_P0_D;
  reg  tlb_6_P0_D;
  reg  tlb_7_P0_D;
  reg  tlb_8_P0_D;
  reg  tlb_9_P0_D;
  reg  tlb_10_P0_D;
  reg  tlb_11_P0_D;
  reg  tlb_12_P0_D;
  reg  tlb_13_P0_D;
  reg  tlb_14_P0_D;
  reg  tlb_15_P0_D;
  wire  _foundTLB_T_666 = tlbHit_15_1 & tlb_15_P0_D;
  wire  foundTLB_1_P0_D = tlbHit_0_1 & tlb_0_P0_D | tlbHit_1_1 & tlb_1_P0_D | tlbHit_2_1 & tlb_2_P0_D | tlbHit_3_1 &
    tlb_3_P0_D | tlbHit_4_1 & tlb_4_P0_D | tlbHit_5_1 & tlb_5_P0_D | tlbHit_6_1 & tlb_6_P0_D | tlbHit_7_1 & tlb_7_P0_D
     | tlbHit_8_1 & tlb_8_P0_D | tlbHit_9_1 & tlb_9_P0_D | tlbHit_10_1 & tlb_10_P0_D | tlbHit_11_1 & tlb_11_P0_D |
    tlbHit_12_1 & tlb_12_P0_D | tlbHit_13_1 & tlb_13_P0_D | tlbHit_14_1 & tlb_14_P0_D | _foundTLB_T_666;
  wire  foundP_1_D = oddPG_1 ? foundTLB_1_P1_D : foundTLB_1_P0_D;
  wire  _GEN_84 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? 1'h0 : ~foundP_1_D;
  wire  pme_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ? 1'h0
     : _GEN_84;
  wire [1:0] _T_626 = _T_135 ? 2'h1 : 2'h0;
  wire [1:0] _T_627 = _T_133 ? 2'h1 : _T_626;
  wire [1:0] _T_628 = _T_131 ? 2'h1 : _T_627;
  wire [1:0] _T_629 = _T_129 ? 2'h0 : _T_628;
  wire [1:0] _T_630 = _T_127 ? 2'h0 : _T_629;
  wire [1:0] _T_631 = _T_125 ? 2'h0 : _T_630;
  wire [1:0] _T_632 = _T_123 ? 2'h3 : _T_631;
  wire [1:0] _T_633 = _T_121 ? 2'h2 : _T_632;
  wire [1:0] _T_634 = _T_119 ? 2'h0 : _T_633;
  wire [1:0] _T_635 = _T_117 ? 2'h0 : _T_634;
  wire [1:0] _T_636 = _T_115 ? 2'h0 : _T_635;
  wire [1:0] _T_637 = _T_113 ? 2'h0 : _T_636;
  wire [1:0] _T_638 = _T_111 ? 2'h0 : _T_637;
  wire [1:0] _T_639 = _T_109 ? 2'h0 : _T_638;
  wire [1:0] _T_640 = _T_107 ? 2'h0 : _T_639;
  wire [1:0] _T_641 = _T_105 ? 2'h0 : _T_640;
  wire [1:0] _T_642 = _T_103 ? 2'h0 : _T_641;
  wire [1:0] _T_643 = _T_101 ? 2'h0 : _T_642;
  wire [1:0] _T_644 = _T_99 ? 2'h0 : _T_643;
  wire [1:0] _T_645 = _T_97 ? 2'h0 : _T_644;
  wire [1:0] _T_646 = _T_95 ? 2'h0 : _T_645;
  wire [1:0] _T_647 = _T_93 ? 2'h0 : _T_646;
  wire [1:0] _T_648 = _T_91 ? 2'h0 : _T_647;
  wire [1:0] _T_649 = _T_89 ? 2'h0 : _T_648;
  wire [1:0] _T_650 = _T_87 ? 2'h0 : _T_649;
  wire [1:0] _T_651 = _T_85 ? 2'h0 : _T_650;
  wire [1:0] _T_652 = _T_83 ? 2'h0 : _T_651;
  wire [1:0] _T_653 = _T_81 ? 2'h0 : _T_652;
  wire [1:0] _T_654 = _T_79 ? 2'h0 : _T_653;
  wire [1:0] _T_655 = _T_77 ? 2'h0 : _T_654;
  wire [1:0] _T_656 = _T_75 ? 2'h0 : _T_655;
  wire [1:0] _T_657 = _T_73 ? 2'h0 : _T_656;
  wire [1:0] _T_658 = _T_71 ? 2'h0 : _T_657;
  wire [1:0] _T_659 = _T_69 ? 2'h0 : _T_658;
  wire [1:0] _T_660 = _T_67 ? 2'h0 : _T_659;
  wire [1:0] _T_661 = _T_65 ? 2'h0 : _T_660;
  wire [1:0] _T_662 = _T_63 ? 2'h0 : _T_661;
  wire [1:0] _T_663 = _T_61 ? 2'h0 : _T_662;
  wire [1:0] _T_664 = _T_59 ? 2'h0 : _T_663;
  wire [1:0] _T_665 = _T_57 ? 2'h0 : _T_664;
  wire [1:0] _T_666 = _T_55 ? 2'h0 : _T_665;
  wire [1:0] _T_667 = _T_53 ? 2'h0 : _T_666;
  wire [1:0] _T_668 = _T_51 ? 2'h0 : _T_667;
  wire [1:0] _T_669 = _T_49 ? 2'h0 : _T_668;
  wire [1:0] _T_670 = _T_47 ? 2'h0 : _T_669;
  wire [1:0] _T_671 = _T_45 ? 2'h0 : _T_670;
  wire [1:0] _T_672 = _T_43 ? 2'h0 : _T_671;
  wire [1:0] _T_673 = _T_41 ? 2'h0 : _T_672;
  wire [1:0] _T_674 = _T_39 ? 2'h0 : _T_673;
  wire [1:0] _T_675 = _T_37 ? 2'h0 : _T_674;
  wire [1:0] c0_2 = _T_35 ? 2'h0 : _T_675;
  wire  _GEN_99 = pme_1 & c0_2[0] & _TLBR_T;
  wire  _GEN_103 = ppi_1 ? 1'h0 : _GEN_99;
  wire  _GEN_109 = invalid_1 ? 1'h0 : _GEN_103;
  wire  _GEN_116 = miss_1 ? 1'h0 : _GEN_109;
  wire  _GEN_133 = crmd_DA ? 1'h0 : _GEN_116;
  wire  _GEN_142 = memALE ? 1'h0 : _GEN_133;
  wire  _GEN_151 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_142;
  wire  _GEN_163 = ID_OK & _GEN_151;
  wire  PME = dStallReg ? 1'h0 : _GEN_163;
  wire  _GEN_23 = invalid ? 1'h0 : ppi;
  wire  _GEN_27 = miss ? 1'h0 : _GEN_23;
  wire  _GEN_38 = crmd_DA ? 1'h0 : _GEN_27;
  wire  _GEN_43 = PC[1:0] != 2'h0 ? 1'h0 : _GEN_38;
  wire  _GEN_51 = ~INT & ~idle & _GEN_43;
  wire  _GEN_58 = dStallReg | iStallReg ? 1'h0 : _GEN_51;
  wire  _GEN_102 = ppi_1 ? _TLBR_T : _GEN_58;
  wire  _GEN_108 = invalid_1 ? _GEN_58 : _GEN_102;
  wire  _GEN_115 = miss_1 ? _GEN_58 : _GEN_108;
  wire  _GEN_132 = crmd_DA ? _GEN_58 : _GEN_115;
  wire  _GEN_141 = memALE ? _GEN_58 : _GEN_132;
  wire  _GEN_150 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? _GEN_58 : _GEN_141;
  wire  _GEN_162 = ID_OK ? _GEN_150 : _GEN_58;
  wire  PPI = dStallReg ? _GEN_58 : _GEN_162;
  wire  _GEN_97 = c0_2[0] & _TLBR_T;
  wire  _GEN_106 = invalid_1 & _GEN_97;
  wire  _GEN_113 = miss_1 ? 1'h0 : _GEN_106;
  wire  _GEN_130 = crmd_DA ? 1'h0 : _GEN_113;
  wire  _GEN_139 = memALE ? 1'h0 : _GEN_130;
  wire  _GEN_148 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_139;
  wire  _GEN_160 = ID_OK & _GEN_148;
  wire  PIS = dStallReg ? 1'h0 : _GEN_160;
  wire  _GEN_26 = miss ? 1'h0 : invalid;
  wire  _GEN_37 = crmd_DA ? 1'h0 : _GEN_26;
  wire  _GEN_42 = PC[1:0] != 2'h0 ? 1'h0 : _GEN_37;
  wire  _GEN_50 = ~INT & ~idle & _GEN_42;
  wire  PIF = dStallReg | iStallReg ? 1'h0 : _GEN_50;
  wire  _GEN_98 = c0_2[0] ? 1'h0 : _TLBR_T;
  wire  _GEN_107 = invalid_1 & _GEN_98;
  wire  _GEN_114 = miss_1 ? 1'h0 : _GEN_107;
  wire  _GEN_131 = crmd_DA ? 1'h0 : _GEN_114;
  wire  _GEN_140 = memALE ? 1'h0 : _GEN_131;
  wire  _GEN_149 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? 1'h0 : _GEN_140;
  wire  _GEN_161 = ID_OK & _GEN_149;
  wire  PIL = dStallReg ? 1'h0 : _GEN_161;
  wire [15:0] _excp_T = {INT,PIL,PIS,PIF,PME,PPI,ADEF,1'h0,excp_lo};
  wire  excp = |_excp_T;
  reg [19:0] tlb_0_P0_PPN;
  reg [1:0] tlb_0_P0_MAT;
  reg [19:0] tlb_0_P1_PPN;
  reg [1:0] tlb_0_P1_MAT;
  reg [19:0] tlb_1_P0_PPN;
  reg [1:0] tlb_1_P0_MAT;
  reg [19:0] tlb_1_P1_PPN;
  reg [1:0] tlb_1_P1_MAT;
  reg [19:0] tlb_2_P0_PPN;
  reg [1:0] tlb_2_P0_MAT;
  reg [19:0] tlb_2_P1_PPN;
  reg [1:0] tlb_2_P1_MAT;
  reg [19:0] tlb_3_P0_PPN;
  reg [1:0] tlb_3_P0_MAT;
  reg [19:0] tlb_3_P1_PPN;
  reg [1:0] tlb_3_P1_MAT;
  reg [19:0] tlb_4_P0_PPN;
  reg [1:0] tlb_4_P0_MAT;
  reg [19:0] tlb_4_P1_PPN;
  reg [1:0] tlb_4_P1_MAT;
  reg [19:0] tlb_5_P0_PPN;
  reg [1:0] tlb_5_P0_MAT;
  reg [19:0] tlb_5_P1_PPN;
  reg [1:0] tlb_5_P1_MAT;
  reg [19:0] tlb_6_P0_PPN;
  reg [1:0] tlb_6_P0_MAT;
  reg [19:0] tlb_6_P1_PPN;
  reg [1:0] tlb_6_P1_MAT;
  reg [19:0] tlb_7_P0_PPN;
  reg [1:0] tlb_7_P0_MAT;
  reg [19:0] tlb_7_P1_PPN;
  reg [1:0] tlb_7_P1_MAT;
  reg [19:0] tlb_8_P0_PPN;
  reg [1:0] tlb_8_P0_MAT;
  reg [19:0] tlb_8_P1_PPN;
  reg [1:0] tlb_8_P1_MAT;
  reg [19:0] tlb_9_P0_PPN;
  reg [1:0] tlb_9_P0_MAT;
  reg [19:0] tlb_9_P1_PPN;
  reg [1:0] tlb_9_P1_MAT;
  reg [19:0] tlb_10_P0_PPN;
  reg [1:0] tlb_10_P0_MAT;
  reg [19:0] tlb_10_P1_PPN;
  reg [1:0] tlb_10_P1_MAT;
  reg [19:0] tlb_11_P0_PPN;
  reg [1:0] tlb_11_P0_MAT;
  reg [19:0] tlb_11_P1_PPN;
  reg [1:0] tlb_11_P1_MAT;
  reg [19:0] tlb_12_P0_PPN;
  reg [1:0] tlb_12_P0_MAT;
  reg [19:0] tlb_12_P1_PPN;
  reg [1:0] tlb_12_P1_MAT;
  reg [19:0] tlb_13_P0_PPN;
  reg [1:0] tlb_13_P0_MAT;
  reg [19:0] tlb_13_P1_PPN;
  reg [1:0] tlb_13_P1_MAT;
  reg [19:0] tlb_14_P0_PPN;
  reg [1:0] tlb_14_P0_MAT;
  reg [19:0] tlb_14_P1_PPN;
  reg [1:0] tlb_14_P1_MAT;
  reg [19:0] tlb_15_P0_PPN;
  reg [1:0] tlb_15_P0_MAT;
  reg [19:0] tlb_15_P1_PPN;
  reg [1:0] tlb_15_P1_MAT;
  wire [31:0] _pa_T_1 = {csrs_27_PSEG,PC[28:0]};
  wire [31:0] _pa_T_3 = {csrs_28_PSEG,PC[28:0]};
  wire [19:0] _foundTLB_T_124 = tlbHit_0 ? tlb_0_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_125 = tlbHit_1 ? tlb_1_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_126 = tlbHit_2 ? tlb_2_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_127 = tlbHit_3 ? tlb_3_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_128 = tlbHit_4 ? tlb_4_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_129 = tlbHit_5 ? tlb_5_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_130 = tlbHit_6 ? tlb_6_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_131 = tlbHit_7 ? tlb_7_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_132 = tlbHit_8 ? tlb_8_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_133 = tlbHit_9 ? tlb_9_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_134 = tlbHit_10 ? tlb_10_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_135 = tlbHit_11 ? tlb_11_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_136 = tlbHit_12 ? tlb_12_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_137 = tlbHit_13 ? tlb_13_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_138 = tlbHit_14 ? tlb_14_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_139 = tlbHit_15 ? tlb_15_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_140 = _foundTLB_T_124 | _foundTLB_T_125;
  wire [19:0] _foundTLB_T_141 = _foundTLB_T_140 | _foundTLB_T_126;
  wire [19:0] _foundTLB_T_142 = _foundTLB_T_141 | _foundTLB_T_127;
  wire [19:0] _foundTLB_T_143 = _foundTLB_T_142 | _foundTLB_T_128;
  wire [19:0] _foundTLB_T_144 = _foundTLB_T_143 | _foundTLB_T_129;
  wire [19:0] _foundTLB_T_145 = _foundTLB_T_144 | _foundTLB_T_130;
  wire [19:0] _foundTLB_T_146 = _foundTLB_T_145 | _foundTLB_T_131;
  wire [19:0] _foundTLB_T_147 = _foundTLB_T_146 | _foundTLB_T_132;
  wire [19:0] _foundTLB_T_148 = _foundTLB_T_147 | _foundTLB_T_133;
  wire [19:0] _foundTLB_T_149 = _foundTLB_T_148 | _foundTLB_T_134;
  wire [19:0] _foundTLB_T_150 = _foundTLB_T_149 | _foundTLB_T_135;
  wire [19:0] _foundTLB_T_151 = _foundTLB_T_150 | _foundTLB_T_136;
  wire [19:0] _foundTLB_T_152 = _foundTLB_T_151 | _foundTLB_T_137;
  wire [19:0] _foundTLB_T_153 = _foundTLB_T_152 | _foundTLB_T_138;
  wire [19:0] foundTLB_P1_PPN = _foundTLB_T_153 | _foundTLB_T_139;
  wire [19:0] _foundTLB_T_279 = tlbHit_0 ? tlb_0_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_280 = tlbHit_1 ? tlb_1_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_281 = tlbHit_2 ? tlb_2_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_282 = tlbHit_3 ? tlb_3_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_283 = tlbHit_4 ? tlb_4_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_284 = tlbHit_5 ? tlb_5_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_285 = tlbHit_6 ? tlb_6_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_286 = tlbHit_7 ? tlb_7_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_287 = tlbHit_8 ? tlb_8_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_288 = tlbHit_9 ? tlb_9_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_289 = tlbHit_10 ? tlb_10_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_290 = tlbHit_11 ? tlb_11_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_291 = tlbHit_12 ? tlb_12_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_292 = tlbHit_13 ? tlb_13_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_293 = tlbHit_14 ? tlb_14_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_294 = tlbHit_15 ? tlb_15_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_295 = _foundTLB_T_279 | _foundTLB_T_280;
  wire [19:0] _foundTLB_T_296 = _foundTLB_T_295 | _foundTLB_T_281;
  wire [19:0] _foundTLB_T_297 = _foundTLB_T_296 | _foundTLB_T_282;
  wire [19:0] _foundTLB_T_298 = _foundTLB_T_297 | _foundTLB_T_283;
  wire [19:0] _foundTLB_T_299 = _foundTLB_T_298 | _foundTLB_T_284;
  wire [19:0] _foundTLB_T_300 = _foundTLB_T_299 | _foundTLB_T_285;
  wire [19:0] _foundTLB_T_301 = _foundTLB_T_300 | _foundTLB_T_286;
  wire [19:0] _foundTLB_T_302 = _foundTLB_T_301 | _foundTLB_T_287;
  wire [19:0] _foundTLB_T_303 = _foundTLB_T_302 | _foundTLB_T_288;
  wire [19:0] _foundTLB_T_304 = _foundTLB_T_303 | _foundTLB_T_289;
  wire [19:0] _foundTLB_T_305 = _foundTLB_T_304 | _foundTLB_T_290;
  wire [19:0] _foundTLB_T_306 = _foundTLB_T_305 | _foundTLB_T_291;
  wire [19:0] _foundTLB_T_307 = _foundTLB_T_306 | _foundTLB_T_292;
  wire [19:0] _foundTLB_T_308 = _foundTLB_T_307 | _foundTLB_T_293;
  wire [19:0] foundTLB_P0_PPN = _foundTLB_T_308 | _foundTLB_T_294;
  wire [19:0] foundP_PPN = oddPG ? foundTLB_P1_PPN : foundTLB_P0_PPN;
  wire [31:0] _pa_T_6 = {foundP_PPN,PC[11:0]};
  wire [21:0] _pa_T_9 = {foundP_PPN[19:9],PC[20:10]};
  wire [31:0] _pa_T_10 = _oddPG_T ? _pa_T_6 : {{10'd0}, _pa_T_9};
  wire [31:0] _GEN_6 = PC[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? _pa_T_3 : _pa_T_10;
  wire [31:0] pa = PC[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3) ?
    _pa_T_1 : _GEN_6;
  wire  _io_inst_req_valid_T_1 = ~dStallReg;
  wire [18:0] _GEN_44 = ~ADEF ? PC[31:13] : csrs_9_VPPN;
  wire [31:0] _GEN_45 = ~IF_OK ? PC : badv_VAddr;
  wire [18:0] _GEN_46 = ~IF_OK ? _GEN_44 : csrs_9_VPPN;
  wire [31:0] _GEN_52 = ~INT & ~idle ? _GEN_45 : badv_VAddr;
  wire [18:0] _GEN_53 = ~INT & ~idle ? _GEN_46 : csrs_9_VPPN;
  wire [31:0] _GEN_59 = dStallReg | iStallReg ? badv_VAddr : _GEN_52;
  wire [18:0] _GEN_60 = dStallReg | iStallReg ? csrs_9_VPPN : _GEN_53;
  wire [2:0] _T_490 = _T_151 ? 3'h2 : 3'h0;
  wire [2:0] _T_491 = _T_149 ? 3'h0 : _T_490;
  wire [2:0] _T_492 = _T_147 ? 3'h2 : _T_491;
  wire [2:0] _T_493 = _T_145 ? 3'h0 : _T_492;
  wire [2:0] _T_494 = _T_143 ? 3'h0 : _T_493;
  wire [2:0] _T_495 = _T_141 ? 3'h0 : _T_494;
  wire [2:0] _T_496 = _T_139 ? 3'h1 : _T_495;
  wire [2:0] _T_497 = _T_137 ? 3'h1 : _T_496;
  wire [2:0] _T_498 = _T_135 ? 3'h0 : _T_497;
  wire [2:0] _T_499 = _T_133 ? 3'h0 : _T_498;
  wire [2:0] _T_500 = _T_131 ? 3'h0 : _T_499;
  wire [2:0] _T_501 = _T_129 ? 3'h1 : _T_500;
  wire [2:0] _T_502 = _T_127 ? 3'h1 : _T_501;
  wire [2:0] _T_503 = _T_125 ? 3'h1 : _T_502;
  wire [2:0] _T_504 = _T_123 ? 3'h7 : _T_503;
  wire [2:0] _T_505 = _T_121 ? 3'h1 : _T_504;
  wire [2:0] _T_506 = _T_119 ? 3'h0 : _T_505;
  wire [2:0] _T_507 = _T_117 ? 3'h0 : _T_506;
  wire [2:0] _T_508 = _T_115 ? 3'h0 : _T_507;
  wire [2:0] _T_509 = _T_113 ? 3'h0 : _T_508;
  wire [2:0] _T_510 = _T_111 ? 3'h0 : _T_509;
  wire [2:0] _T_511 = _T_109 ? 3'h0 : _T_510;
  wire [2:0] _T_512 = _T_107 ? 3'h0 : _T_511;
  wire [2:0] _T_513 = _T_105 ? 3'h0 : _T_512;
  wire [2:0] _T_514 = _T_103 ? 3'h0 : _T_513;
  wire [2:0] _T_515 = _T_101 ? 3'h0 : _T_514;
  wire [2:0] _T_516 = _T_99 ? 3'h3 : _T_515;
  wire [2:0] _T_517 = _T_97 ? 3'h0 : _T_516;
  wire [2:0] _T_518 = _T_95 ? 3'h0 : _T_517;
  wire [2:0] _T_519 = _T_93 ? 3'h0 : _T_518;
  wire [2:0] _T_520 = _T_91 ? 3'h0 : _T_519;
  wire [2:0] _T_521 = _T_89 ? 3'h0 : _T_520;
  wire [2:0] _T_522 = _T_87 ? 3'h0 : _T_521;
  wire [2:0] _T_523 = _T_85 ? 3'h0 : _T_522;
  wire [2:0] _T_524 = _T_83 ? 3'h0 : _T_523;
  wire [2:0] _T_525 = _T_81 ? 3'h0 : _T_524;
  wire [2:0] _T_526 = _T_79 ? 3'h0 : _T_525;
  wire [2:0] _T_527 = _T_77 ? 3'h0 : _T_526;
  wire [2:0] _T_528 = _T_75 ? 3'h0 : _T_527;
  wire [2:0] _T_529 = _T_73 ? 3'h0 : _T_528;
  wire [2:0] _T_530 = _T_71 ? 3'h0 : _T_529;
  wire [2:0] _T_531 = _T_69 ? 3'h0 : _T_530;
  wire [2:0] _T_532 = _T_67 ? 3'h0 : _T_531;
  wire [2:0] _T_533 = _T_65 ? 3'h0 : _T_532;
  wire [2:0] _T_534 = _T_63 ? 3'h0 : _T_533;
  wire [2:0] _T_535 = _T_61 ? 3'h0 : _T_534;
  wire [2:0] _T_536 = _T_59 ? 3'h0 : _T_535;
  wire [2:0] _T_537 = _T_57 ? 3'h0 : _T_536;
  wire [2:0] _T_538 = _T_55 ? 3'h0 : _T_537;
  wire [2:0] _T_539 = _T_53 ? 3'h0 : _T_538;
  wire [2:0] _T_540 = _T_51 ? 3'h0 : _T_539;
  wire [2:0] _T_541 = _T_49 ? 3'h0 : _T_540;
  wire [2:0] _T_542 = _T_47 ? 3'h0 : _T_541;
  wire [2:0] _T_543 = _T_45 ? 3'h0 : _T_542;
  wire [2:0] _T_544 = _T_43 ? 3'h0 : _T_543;
  wire [2:0] _T_545 = _T_41 ? 3'h0 : _T_544;
  wire [2:0] _T_546 = _T_39 ? 3'h5 : _T_545;
  wire [2:0] _T_547 = _T_37 ? 3'h6 : _T_546;
  wire [2:0] c0_0 = _T_35 ? 3'h4 : _T_547;
  wire [1:0] _T_554 = _T_151 ? 2'h1 : 2'h0;
  wire [1:0] _T_555 = _T_149 ? 2'h0 : _T_554;
  wire [1:0] _T_556 = _T_147 ? 2'h2 : _T_555;
  wire [1:0] _T_557 = _T_145 ? 2'h0 : _T_556;
  wire [1:0] _T_558 = _T_143 ? 2'h0 : _T_557;
  wire [1:0] _T_559 = _T_141 ? 2'h0 : _T_558;
  wire [1:0] _T_560 = _T_139 ? 2'h2 : _T_559;
  wire [1:0] _T_561 = _T_137 ? 2'h2 : _T_560;
  wire [1:0] _T_562 = _T_135 ? 2'h0 : _T_561;
  wire [1:0] _T_563 = _T_133 ? 2'h0 : _T_562;
  wire [1:0] _T_564 = _T_131 ? 2'h0 : _T_563;
  wire [1:0] _T_565 = _T_129 ? 2'h2 : _T_564;
  wire [1:0] _T_566 = _T_127 ? 2'h2 : _T_565;
  wire [1:0] _T_567 = _T_125 ? 2'h2 : _T_566;
  wire [1:0] _T_568 = _T_123 ? 2'h2 : _T_567;
  wire [1:0] _T_569 = _T_121 ? 2'h2 : _T_568;
  wire [1:0] _T_570 = _T_119 ? 2'h2 : _T_569;
  wire [1:0] _T_571 = _T_117 ? 2'h2 : _T_570;
  wire [1:0] _T_572 = _T_115 ? 2'h0 : _T_571;
  wire [1:0] _T_573 = _T_113 ? 2'h0 : _T_572;
  wire [1:0] _T_574 = _T_111 ? 2'h0 : _T_573;
  wire [1:0] _T_575 = _T_109 ? 2'h0 : _T_574;
  wire [1:0] _T_576 = _T_107 ? 2'h0 : _T_575;
  wire [1:0] _T_577 = _T_105 ? 2'h0 : _T_576;
  wire [1:0] _T_578 = _T_103 ? 2'h0 : _T_577;
  wire [1:0] _T_579 = _T_101 ? 2'h0 : _T_578;
  wire [1:0] _T_580 = _T_99 ? 2'h2 : _T_579;
  wire [1:0] _T_581 = _T_97 ? 2'h2 : _T_580;
  wire [1:0] _T_582 = _T_95 ? 2'h2 : _T_581;
  wire [1:0] _T_583 = _T_93 ? 2'h2 : _T_582;
  wire [1:0] _T_584 = _T_91 ? 2'h2 : _T_583;
  wire [1:0] _T_585 = _T_89 ? 2'h2 : _T_584;
  wire [1:0] _T_586 = _T_87 ? 2'h2 : _T_585;
  wire [1:0] _T_587 = _T_85 ? 2'h2 : _T_586;
  wire [1:0] _T_588 = _T_83 ? 2'h2 : _T_587;
  wire [1:0] _T_589 = _T_81 ? 2'h2 : _T_588;
  wire [1:0] _T_590 = _T_79 ? 2'h0 : _T_589;
  wire [1:0] _T_591 = _T_77 ? 2'h0 : _T_590;
  wire [1:0] _T_592 = _T_75 ? 2'h2 : _T_591;
  wire [1:0] _T_593 = _T_73 ? 2'h2 : _T_592;
  wire [1:0] _T_594 = _T_71 ? 2'h2 : _T_593;
  wire [1:0] _T_595 = _T_69 ? 2'h2 : _T_594;
  wire [1:0] _T_596 = _T_67 ? 2'h2 : _T_595;
  wire [1:0] _T_597 = _T_65 ? 2'h2 : _T_596;
  wire [1:0] _T_598 = _T_63 ? 2'h2 : _T_597;
  wire [1:0] _T_599 = _T_61 ? 2'h2 : _T_598;
  wire [1:0] _T_600 = _T_59 ? 2'h2 : _T_599;
  wire [1:0] _T_601 = _T_57 ? 2'h2 : _T_600;
  wire [1:0] _T_602 = _T_55 ? 2'h2 : _T_601;
  wire [1:0] _T_603 = _T_53 ? 2'h2 : _T_602;
  wire [1:0] _T_604 = _T_51 ? 2'h2 : _T_603;
  wire [1:0] _T_605 = _T_49 ? 2'h2 : _T_604;
  wire [1:0] _T_606 = _T_47 ? 2'h2 : _T_605;
  wire [1:0] _T_607 = _T_45 ? 2'h2 : _T_606;
  wire [1:0] _T_608 = _T_43 ? 2'h2 : _T_607;
  wire [1:0] _T_609 = _T_41 ? 2'h2 : _T_608;
  wire [1:0] _T_610 = _T_39 ? 2'h2 : _T_609;
  wire [1:0] _T_611 = _T_37 ? 2'h2 : _T_610;
  wire [1:0] c0_1 = _T_35 ? 2'h3 : _T_611;
  wire  _T_1022 = _T_111 ? 1'h0 : _T_113;
  wire  _T_1023 = _T_109 ? 1'h0 : _T_1022;
  wire  _T_1024 = _T_107 ? 1'h0 : _T_1023;
  wire  _T_1025 = _T_105 ? 1'h0 : _T_1024;
  wire  _T_1026 = _T_103 ? 1'h0 : _T_1025;
  wire  _T_1027 = _T_101 ? 1'h0 : _T_1026;
  wire  _T_1028 = _T_99 ? 1'h0 : _T_1027;
  wire  _T_1029 = _T_97 ? 1'h0 : _T_1028;
  wire  _T_1030 = _T_95 ? 1'h0 : _T_1029;
  wire  _T_1031 = _T_93 ? 1'h0 : _T_1030;
  wire  _T_1032 = _T_91 ? 1'h0 : _T_1031;
  wire  _T_1033 = _T_89 ? 1'h0 : _T_1032;
  wire  _T_1034 = _T_87 ? 1'h0 : _T_1033;
  wire  _T_1035 = _T_85 ? 1'h0 : _T_1034;
  wire  _T_1036 = _T_83 ? 1'h0 : _T_1035;
  wire  _T_1037 = _T_81 ? 1'h0 : _T_1036;
  wire  _T_1038 = _T_79 ? 1'h0 : _T_1037;
  wire  _T_1039 = _T_77 ? 1'h0 : _T_1038;
  wire  _T_1040 = _T_75 ? 1'h0 : _T_1039;
  wire  _T_1041 = _T_73 ? 1'h0 : _T_1040;
  wire  _T_1042 = _T_71 ? 1'h0 : _T_1041;
  wire  _T_1043 = _T_69 ? 1'h0 : _T_1042;
  wire  _T_1044 = _T_67 ? 1'h0 : _T_1043;
  wire  _T_1045 = _T_65 ? 1'h0 : _T_1044;
  wire  _T_1046 = _T_63 ? 1'h0 : _T_1045;
  wire  _T_1047 = _T_61 ? 1'h0 : _T_1046;
  wire  _T_1048 = _T_59 ? 1'h0 : _T_1047;
  wire  _T_1049 = _T_57 ? 1'h0 : _T_1048;
  wire  _T_1050 = _T_55 ? 1'h0 : _T_1049;
  wire  _T_1051 = _T_53 ? 1'h0 : _T_1050;
  wire  _T_1052 = _T_51 ? 1'h0 : _T_1051;
  wire  _T_1053 = _T_49 ? 1'h0 : _T_1052;
  wire  _T_1054 = _T_47 ? 1'h0 : _T_1053;
  wire  _T_1055 = _T_45 ? 1'h0 : _T_1054;
  wire  _T_1056 = _T_43 ? 1'h0 : _T_1055;
  wire  _T_1057 = _T_41 ? 1'h0 : _T_1056;
  wire  _T_1058 = _T_39 ? 1'h0 : _T_1057;
  wire  _T_1059 = _T_37 ? 1'h0 : _T_1058;
  wire  c0_8 = _T_35 ? 1'h0 : _T_1059;
  wire  _T_1085 = _T_113 ? 1'h0 : _T_115;
  wire  _T_1086 = _T_111 ? 1'h0 : _T_1085;
  wire  _T_1087 = _T_109 ? 1'h0 : _T_1086;
  wire  _T_1088 = _T_107 ? 1'h0 : _T_1087;
  wire  _T_1089 = _T_105 ? 1'h0 : _T_1088;
  wire  _T_1090 = _T_103 ? 1'h0 : _T_1089;
  wire  _T_1091 = _T_101 ? 1'h0 : _T_1090;
  wire  _T_1092 = _T_99 ? 1'h0 : _T_1091;
  wire  _T_1093 = _T_97 ? 1'h0 : _T_1092;
  wire  _T_1094 = _T_95 ? 1'h0 : _T_1093;
  wire  _T_1095 = _T_93 ? 1'h0 : _T_1094;
  wire  _T_1096 = _T_91 ? 1'h0 : _T_1095;
  wire  _T_1097 = _T_89 ? 1'h0 : _T_1096;
  wire  _T_1098 = _T_87 ? 1'h0 : _T_1097;
  wire  _T_1099 = _T_85 ? 1'h0 : _T_1098;
  wire  _T_1100 = _T_83 ? 1'h0 : _T_1099;
  wire  _T_1101 = _T_81 ? 1'h0 : _T_1100;
  wire  _T_1102 = _T_79 ? 1'h0 : _T_1101;
  wire  _T_1103 = _T_77 ? 1'h0 : _T_1102;
  wire  _T_1104 = _T_75 ? 1'h0 : _T_1103;
  wire  _T_1105 = _T_73 ? 1'h0 : _T_1104;
  wire  _T_1106 = _T_71 ? 1'h0 : _T_1105;
  wire  _T_1107 = _T_69 ? 1'h0 : _T_1106;
  wire  _T_1108 = _T_67 ? 1'h0 : _T_1107;
  wire  _T_1109 = _T_65 ? 1'h0 : _T_1108;
  wire  _T_1110 = _T_63 ? 1'h0 : _T_1109;
  wire  _T_1111 = _T_61 ? 1'h0 : _T_1110;
  wire  _T_1112 = _T_59 ? 1'h0 : _T_1111;
  wire  _T_1113 = _T_57 ? 1'h0 : _T_1112;
  wire  _T_1114 = _T_55 ? 1'h0 : _T_1113;
  wire  _T_1115 = _T_53 ? 1'h0 : _T_1114;
  wire  _T_1116 = _T_51 ? 1'h0 : _T_1115;
  wire  _T_1117 = _T_49 ? 1'h0 : _T_1116;
  wire  _T_1118 = _T_47 ? 1'h0 : _T_1117;
  wire  _T_1119 = _T_45 ? 1'h0 : _T_1118;
  wire  _T_1120 = _T_43 ? 1'h0 : _T_1119;
  wire  _T_1121 = _T_41 ? 1'h0 : _T_1120;
  wire  _T_1122 = _T_39 ? 1'h0 : _T_1121;
  wire  _T_1123 = _T_37 ? 1'h0 : _T_1122;
  wire  c0_9 = _T_35 ? 1'h0 : _T_1123;
  wire [31:0] _pa_T_12 = {csrs_27_PSEG,EXVA[28:0]};
  wire [31:0] _pa_T_14 = {csrs_28_PSEG,EXVA[28:0]};
  wire [19:0] _foundTLB_T_589 = tlbHit_0_1 ? tlb_0_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_590 = tlbHit_1_1 ? tlb_1_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_591 = tlbHit_2_1 ? tlb_2_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_592 = tlbHit_3_1 ? tlb_3_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_593 = tlbHit_4_1 ? tlb_4_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_594 = tlbHit_5_1 ? tlb_5_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_595 = tlbHit_6_1 ? tlb_6_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_596 = tlbHit_7_1 ? tlb_7_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_597 = tlbHit_8_1 ? tlb_8_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_598 = tlbHit_9_1 ? tlb_9_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_599 = tlbHit_10_1 ? tlb_10_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_600 = tlbHit_11_1 ? tlb_11_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_601 = tlbHit_12_1 ? tlb_12_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_602 = tlbHit_13_1 ? tlb_13_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_603 = tlbHit_14_1 ? tlb_14_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_604 = tlbHit_15_1 ? tlb_15_P1_PPN : 20'h0;
  wire [19:0] _foundTLB_T_605 = _foundTLB_T_589 | _foundTLB_T_590;
  wire [19:0] _foundTLB_T_606 = _foundTLB_T_605 | _foundTLB_T_591;
  wire [19:0] _foundTLB_T_607 = _foundTLB_T_606 | _foundTLB_T_592;
  wire [19:0] _foundTLB_T_608 = _foundTLB_T_607 | _foundTLB_T_593;
  wire [19:0] _foundTLB_T_609 = _foundTLB_T_608 | _foundTLB_T_594;
  wire [19:0] _foundTLB_T_610 = _foundTLB_T_609 | _foundTLB_T_595;
  wire [19:0] _foundTLB_T_611 = _foundTLB_T_610 | _foundTLB_T_596;
  wire [19:0] _foundTLB_T_612 = _foundTLB_T_611 | _foundTLB_T_597;
  wire [19:0] _foundTLB_T_613 = _foundTLB_T_612 | _foundTLB_T_598;
  wire [19:0] _foundTLB_T_614 = _foundTLB_T_613 | _foundTLB_T_599;
  wire [19:0] _foundTLB_T_615 = _foundTLB_T_614 | _foundTLB_T_600;
  wire [19:0] _foundTLB_T_616 = _foundTLB_T_615 | _foundTLB_T_601;
  wire [19:0] _foundTLB_T_617 = _foundTLB_T_616 | _foundTLB_T_602;
  wire [19:0] _foundTLB_T_618 = _foundTLB_T_617 | _foundTLB_T_603;
  wire [19:0] foundTLB_1_P1_PPN = _foundTLB_T_618 | _foundTLB_T_604;
  wire [19:0] _foundTLB_T_744 = tlbHit_0_1 ? tlb_0_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_745 = tlbHit_1_1 ? tlb_1_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_746 = tlbHit_2_1 ? tlb_2_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_747 = tlbHit_3_1 ? tlb_3_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_748 = tlbHit_4_1 ? tlb_4_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_749 = tlbHit_5_1 ? tlb_5_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_750 = tlbHit_6_1 ? tlb_6_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_751 = tlbHit_7_1 ? tlb_7_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_752 = tlbHit_8_1 ? tlb_8_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_753 = tlbHit_9_1 ? tlb_9_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_754 = tlbHit_10_1 ? tlb_10_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_755 = tlbHit_11_1 ? tlb_11_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_756 = tlbHit_12_1 ? tlb_12_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_757 = tlbHit_13_1 ? tlb_13_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_758 = tlbHit_14_1 ? tlb_14_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_759 = tlbHit_15_1 ? tlb_15_P0_PPN : 20'h0;
  wire [19:0] _foundTLB_T_760 = _foundTLB_T_744 | _foundTLB_T_745;
  wire [19:0] _foundTLB_T_761 = _foundTLB_T_760 | _foundTLB_T_746;
  wire [19:0] _foundTLB_T_762 = _foundTLB_T_761 | _foundTLB_T_747;
  wire [19:0] _foundTLB_T_763 = _foundTLB_T_762 | _foundTLB_T_748;
  wire [19:0] _foundTLB_T_764 = _foundTLB_T_763 | _foundTLB_T_749;
  wire [19:0] _foundTLB_T_765 = _foundTLB_T_764 | _foundTLB_T_750;
  wire [19:0] _foundTLB_T_766 = _foundTLB_T_765 | _foundTLB_T_751;
  wire [19:0] _foundTLB_T_767 = _foundTLB_T_766 | _foundTLB_T_752;
  wire [19:0] _foundTLB_T_768 = _foundTLB_T_767 | _foundTLB_T_753;
  wire [19:0] _foundTLB_T_769 = _foundTLB_T_768 | _foundTLB_T_754;
  wire [19:0] _foundTLB_T_770 = _foundTLB_T_769 | _foundTLB_T_755;
  wire [19:0] _foundTLB_T_771 = _foundTLB_T_770 | _foundTLB_T_756;
  wire [19:0] _foundTLB_T_772 = _foundTLB_T_771 | _foundTLB_T_757;
  wire [19:0] _foundTLB_T_773 = _foundTLB_T_772 | _foundTLB_T_758;
  wire [19:0] foundTLB_1_P0_PPN = _foundTLB_T_773 | _foundTLB_T_759;
  wire [19:0] foundP_1_PPN = oddPG_1 ? foundTLB_1_P1_PPN : foundTLB_1_P0_PPN;
  wire [31:0] _pa_T_17 = {foundP_1_PPN,EXVA[11:0]};
  wire [21:0] _pa_T_20 = {foundP_1_PPN[19:9],EXVA[20:10]};
  wire [31:0] _pa_T_21 = _oddPG_T_3 ? _pa_T_17 : {{10'd0}, _pa_T_20};
  wire [31:0] _GEN_78 = EXVA[31:29] == csrs_28_VSEG & (csrs_28_PLV0 & _T_12 | csrs_28_PLV3 & _T_14) ? _pa_T_14 :
    _pa_T_21;
  wire [31:0] pa_1 = EXVA[31:29] == csrs_27_VSEG & (csrs_27_PLV0 & crmd_PLV == 2'h0 | csrs_27_PLV3 & crmd_PLV == 2'h3)
     ? _pa_T_12 : _GEN_78;
  wire [3:0] _GEN_93 = 2'h1 == c0_3[2:1] ? 4'h3 : 4'h1;
  wire [3:0] _GEN_94 = 2'h2 == c0_3[2:1] ? 4'hf : _GEN_93;
  wire [3:0] _GEN_95 = 2'h3 == c0_3[2:1] ? 4'h0 : _GEN_94;
  wire [6:0] _GEN_8 = {{3'd0}, _GEN_95};
  wire [6:0] memMask = _GEN_8 << aluOut[1:0];
  wire  _GEN_100 = pme_1 & c0_2[0] ? c0_12 : 1'h1;
  wire  _GEN_104 = ppi_1 ? c0_12 : _GEN_100;
  wire  _GEN_110 = invalid_1 ? c0_12 : _GEN_104;
  wire  _GEN_117 = miss_1 ? c0_12 : _GEN_110;
  wire  _GEN_127 = crmd_DA | _GEN_117;
  wire  _GEN_136 = memALE ? c0_12 : _GEN_127;
  wire  _GEN_144 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 | _GEN_136;
  wire  _GEN_156 = ID_OK & _GEN_144;
  wire  mem_OK = dStallReg | _GEN_156;
  wire  _GEN_101 = pme_1 & c0_2[0] & c0_12;
  wire  _GEN_105 = ppi_1 ? c0_12 : _GEN_101;
  wire  _GEN_111 = invalid_1 ? c0_12 : _GEN_105;
  wire  _GEN_118 = miss_1 ? c0_12 : _GEN_111;
  wire  _GEN_134 = crmd_DA ? c0_12 : _GEN_118;
  wire  _GEN_143 = memALE ? c0_12 : _GEN_134;
  wire  _GEN_152 = c0_3 == 3'h7 | c0_11 & d[4:3] != 2'h2 ? c0_12 : _GEN_143;
  wire  _GEN_164 = ID_OK ? _GEN_152 : c0_12;
  wire  preldNop = dStallReg ? c0_12 : _GEN_164;
  wire  _io_data_req_bits_wen_T_1 = c0_2 == 2'h3;
  wire [6:0] _io_data_req_bits_wen_T_4 = c0_2 == 2'h1 | c0_2 == 2'h3 & csrs_25_ROLLB ? memMask : 7'h0;
  wire [4:0] _io_data_req_bits_wdata_T_1 = {aluOut[1:0], 3'h0};
  wire [62:0] _GEN_12 = {{31'd0}, rkd};
  wire [62:0] _io_data_req_bits_wdata_T_2 = _GEN_12 << _io_data_req_bits_wdata_T_1;
  wire [31:0] shiftData = io_data_resp_bits >> _io_data_req_bits_wdata_T_1;
  wire  _extendData_T = c0_3 == 3'h0;
  wire [23:0] _extendData_T_3 = shiftData[7] ? 24'hffffff : 24'h0;
  wire [31:0] _extendData_T_5 = {_extendData_T_3,shiftData[7:0]};
  wire  _extendData_T_6 = c0_3 == 3'h1;
  wire [31:0] _extendData_T_8 = {24'h0,shiftData[7:0]};
  wire  _extendData_T_9 = c0_3 == 3'h2;
  wire [15:0] _extendData_T_12 = shiftData[15] ? 16'hffff : 16'h0;
  wire [31:0] _extendData_T_14 = {_extendData_T_12,shiftData[15:0]};
  wire  _extendData_T_15 = c0_3 == 3'h3;
  wire [31:0] _extendData_T_17 = {16'h0,shiftData[15:0]};
  wire  _extendData_T_18 = c0_3 == 3'h4;
  wire [31:0] _extendData_T_19 = _extendData_T ? _extendData_T_5 : 32'h0;
  wire [31:0] _extendData_T_20 = _extendData_T_6 ? _extendData_T_8 : 32'h0;
  wire [31:0] _extendData_T_21 = _extendData_T_9 ? _extendData_T_14 : 32'h0;
  wire [31:0] _extendData_T_22 = _extendData_T_15 ? _extendData_T_17 : 32'h0;
  wire [31:0] _extendData_T_23 = _extendData_T_18 ? shiftData : 32'h0;
  wire [31:0] _extendData_T_24 = _extendData_T_19 | _extendData_T_20;
  wire [31:0] _extendData_T_25 = _extendData_T_24 | _extendData_T_21;
  wire [31:0] _extendData_T_26 = _extendData_T_25 | _extendData_T_22;
  wire [31:0] extendData = _extendData_T_26 | _extendData_T_23;
  wire [18:0] _GEN_153 = ~ALE ? aluOut[31:13] : _GEN_60;
  wire [31:0] _GEN_154 = ~mem_OK ? aluOut : _GEN_59;
  wire [18:0] _GEN_155 = ~mem_OK ? _GEN_153 : _GEN_60;
  wire [31:0] _GEN_165 = ID_OK ? _GEN_154 : _GEN_59;
  wire [18:0] _GEN_166 = ID_OK ? _GEN_155 : _GEN_60;
  wire [31:0] _GEN_176 = dStallReg ? _GEN_59 : _GEN_165;
  wire [18:0] _GEN_177 = dStallReg ? _GEN_60 : _GEN_166;
  wire  dStall = ~io_data_resp_valid & (io_data_req_valid | dStallReg);
  wire  _T_1355 = ~dStall;
  wire  _GEN_178 = c0_2 == 2'h2 & mem_OK & ~dStall | csrs_25_ROLLB;
  wire  _GEN_179 = _io_data_req_bits_wen_T_1 & mem_OK & _T_1355 ? 1'h0 : _GEN_178;
  wire  _csrRD_T = 14'h0 == inst[23:10];
  wire [8:0] _csrRD_T_1 = {crmd_DATM,crmd_DATF,crmd_PG,crmd_DA,crmd_IE,crmd_PLV};
  wire  _csrRD_T_2 = 14'h1 == inst[23:10];
  wire [2:0] _csrRD_T_3 = {csrs_1_PIE,csrs_1_PPLV};
  wire  _csrRD_T_4 = 14'h2 == inst[23:10];
  wire  _csrRD_T_5 = 14'h4 == inst[23:10];
  wire  _csrRD_T_6 = 14'h5 == inst[23:10];
  wire [7:0] csrRD_lo_1 = {csrs_4_IS_7,csrs_4_IS_6,csrs_4_IS_5,csrs_4_IS_4,csrs_4_IS_3,csrs_4_IS_2,csrs_4_IS_1,
    csrs_4_IS_0};
  wire [30:0] _csrRD_T_7 = {9'h0,csrs_4_Ecode,3'h0,csrs_4_IS_12,csrs_4_IS_11,1'h0,csrs_4_IS_9,csrs_4_IS_8,csrRD_lo_1};
  wire  _csrRD_T_8 = 14'h6 == inst[23:10];
  wire  _csrRD_T_9 = 14'h7 == inst[23:10];
  wire  _csrRD_T_10 = 14'hc == inst[23:10];
  wire [31:0] _csrRD_T_11 = {csrs_7_VA,6'h0};
  wire  _csrRD_T_12 = 14'h10 == inst[23:10];
  wire [31:0] _csrRD_T_13 = {csrs_8_NE,1'h0,csrs_8_PS,20'h0,csrs_8_Index};
  wire  _csrRD_T_14 = 14'h11 == inst[23:10];
  wire  _csrRD_T_16 = 14'h12 == inst[23:10];
  wire [31:0] _csrRD_T_17 = {csrs_10_PPN,1'h0,csrs_10_G,csrs_10_MAT,csrs_10_PLV,csrs_10_D,csrs_10_V};
  wire  _csrRD_T_18 = 14'h13 == inst[23:10];
  wire [31:0] _csrRD_T_19 = {csrs_11_PPN,1'h0,csrs_11_G,csrs_11_MAT,csrs_11_PLV,csrs_11_D,csrs_11_V};
  wire  _csrRD_T_20 = 14'h18 == inst[23:10];
  wire [23:0] _csrRD_T_21 = {14'h280,asid_ASID};
  wire  _csrRD_T_22 = 14'h19 == inst[23:10];
  wire [31:0] _csrRD_T_23 = {csrs_13_Base,12'h0};
  wire  _csrRD_T_24 = 14'h1a == inst[23:10];
  wire [31:0] _csrRD_T_25 = {csrs_14_Base,12'h0};
  wire  _csrRD_T_26 = 14'h1b == inst[23:10];
  wire [31:0] _csrRD_T_30 = badv_VAddr[31] ? _csrRD_T_25 : _csrRD_T_23;
  wire  _csrRD_T_32 = 14'h30 == inst[23:10];
  wire  _csrRD_T_33 = 14'h31 == inst[23:10];
  wire  _csrRD_T_34 = 14'h32 == inst[23:10];
  wire  _csrRD_T_35 = 14'h33 == inst[23:10];
  wire  _csrRD_T_36 = 14'h40 == inst[23:10];
  wire  _csrRD_T_37 = 14'h41 == inst[23:10];
  wire [31:0] _csrRD_T_38 = {csrs_22_InitVal,csrs_22_Periodic,csrs_22_En};
  wire  _csrRD_T_39 = 14'h42 == inst[23:10];
  wire  _csrRD_T_40 = 14'h44 == inst[23:10];
  wire  _csrRD_T_41 = 14'h60 == inst[23:10];
  wire [2:0] _csrRD_T_42 = {csrs_25_KLO,1'h0,csrs_25_ROLLB};
  wire  _csrRD_T_43 = 14'h88 == inst[23:10];
  wire [31:0] _csrRD_T_44 = {csrs_26_PA,6'h0};
  wire  _csrRD_T_45 = 14'h180 == inst[23:10];
  wire [31:0] _csrRD_T_46 = {csrs_27_VSEG,1'h0,csrs_27_PSEG,19'h0,csrs_27_MAT,csrs_27_PLV3,2'h0,csrs_27_PLV0};
  wire  _csrRD_T_47 = 14'h181 == inst[23:10];
  wire [31:0] _csrRD_T_48 = {csrs_28_VSEG,1'h0,csrs_28_PSEG,19'h0,csrs_28_MAT,csrs_28_PLV3,2'h0,csrs_28_PLV0};
  wire [8:0] _csrRD_T_49 = _csrRD_T ? _csrRD_T_1 : 9'h0;
  wire [2:0] _csrRD_T_50 = _csrRD_T_2 ? _csrRD_T_3 : 3'h0;
  wire  _csrRD_T_51 = _csrRD_T_4 & csrs_2_FPE;
  wire [12:0] _csrRD_T_52 = _csrRD_T_5 ? csrs_3_LIE : 13'h0;
  wire [30:0] _csrRD_T_53 = _csrRD_T_6 ? _csrRD_T_7 : 31'h0;
  wire [31:0] _csrRD_T_54 = _csrRD_T_8 ? csrs_5_PC : 32'h0;
  wire [31:0] _csrRD_T_55 = _csrRD_T_9 ? badv_VAddr : 32'h0;
  wire [31:0] _csrRD_T_56 = _csrRD_T_10 ? _csrRD_T_11 : 32'h0;
  wire [31:0] _csrRD_T_57 = _csrRD_T_12 ? _csrRD_T_13 : 32'h0;
  wire [31:0] _csrRD_T_58 = _csrRD_T_14 ? _EXVA_T_2 : 32'h0;
  wire [31:0] _csrRD_T_59 = _csrRD_T_16 ? _csrRD_T_17 : 32'h0;
  wire [31:0] _csrRD_T_60 = _csrRD_T_18 ? _csrRD_T_19 : 32'h0;
  wire [23:0] _csrRD_T_61 = _csrRD_T_20 ? _csrRD_T_21 : 24'h0;
  wire [31:0] _csrRD_T_62 = _csrRD_T_22 ? _csrRD_T_23 : 32'h0;
  wire [31:0] _csrRD_T_63 = _csrRD_T_24 ? _csrRD_T_25 : 32'h0;
  wire [31:0] _csrRD_T_64 = _csrRD_T_26 ? _csrRD_T_30 : 32'h0;
  wire [31:0] _csrRD_T_66 = _csrRD_T_32 ? csrs_17_Data : 32'h0;
  wire [31:0] _csrRD_T_67 = _csrRD_T_33 ? csrs_18_Data : 32'h0;
  wire [31:0] _csrRD_T_68 = _csrRD_T_34 ? csrs_19_Data : 32'h0;
  wire [31:0] _csrRD_T_69 = _csrRD_T_35 ? csrs_20_Data : 32'h0;
  wire [31:0] _csrRD_T_70 = _csrRD_T_36 ? csrs_21_TID : 32'h0;
  wire [31:0] _csrRD_T_71 = _csrRD_T_37 ? _csrRD_T_38 : 32'h0;
  wire [31:0] _csrRD_T_72 = _csrRD_T_39 ? csrs_23_TimeVal : 32'h0;
  wire [2:0] _csrRD_T_74 = _csrRD_T_41 ? _csrRD_T_42 : 3'h0;
  wire [31:0] _csrRD_T_75 = _csrRD_T_43 ? _csrRD_T_44 : 32'h0;
  wire [31:0] _csrRD_T_76 = _csrRD_T_45 ? _csrRD_T_46 : 32'h0;
  wire [31:0] _csrRD_T_77 = _csrRD_T_47 ? _csrRD_T_48 : 32'h0;
  wire [8:0] _GEN_2359 = {{6'd0}, _csrRD_T_50};
  wire [8:0] _csrRD_T_78 = _csrRD_T_49 | _GEN_2359;
  wire [8:0] _GEN_2360 = {{8'd0}, _csrRD_T_51};
  wire [8:0] _csrRD_T_79 = _csrRD_T_78 | _GEN_2360;
  wire [12:0] _GEN_2361 = {{4'd0}, _csrRD_T_79};
  wire [12:0] _csrRD_T_80 = _GEN_2361 | _csrRD_T_52;
  wire [30:0] _GEN_2362 = {{18'd0}, _csrRD_T_80};
  wire [30:0] _csrRD_T_81 = _GEN_2362 | _csrRD_T_53;
  wire [31:0] _GEN_2363 = {{1'd0}, _csrRD_T_81};
  wire [31:0] _csrRD_T_82 = _GEN_2363 | _csrRD_T_54;
  wire [31:0] _csrRD_T_83 = _csrRD_T_82 | _csrRD_T_55;
  wire [31:0] _csrRD_T_84 = _csrRD_T_83 | _csrRD_T_56;
  wire [31:0] _csrRD_T_85 = _csrRD_T_84 | _csrRD_T_57;
  wire [31:0] _csrRD_T_86 = _csrRD_T_85 | _csrRD_T_58;
  wire [31:0] _csrRD_T_87 = _csrRD_T_86 | _csrRD_T_59;
  wire [31:0] _csrRD_T_88 = _csrRD_T_87 | _csrRD_T_60;
  wire [31:0] _GEN_2364 = {{8'd0}, _csrRD_T_61};
  wire [31:0] _csrRD_T_89 = _csrRD_T_88 | _GEN_2364;
  wire [31:0] _csrRD_T_90 = _csrRD_T_89 | _csrRD_T_62;
  wire [31:0] _csrRD_T_91 = _csrRD_T_90 | _csrRD_T_63;
  wire [31:0] _csrRD_T_92 = _csrRD_T_91 | _csrRD_T_64;
  wire [31:0] _csrRD_T_94 = _csrRD_T_92 | _csrRD_T_66;
  wire [31:0] _csrRD_T_95 = _csrRD_T_94 | _csrRD_T_67;
  wire [31:0] _csrRD_T_96 = _csrRD_T_95 | _csrRD_T_68;
  wire [31:0] _csrRD_T_97 = _csrRD_T_96 | _csrRD_T_69;
  wire [31:0] _csrRD_T_98 = _csrRD_T_97 | _csrRD_T_70;
  wire [31:0] _csrRD_T_99 = _csrRD_T_98 | _csrRD_T_71;
  wire [31:0] _csrRD_T_100 = _csrRD_T_99 | _csrRD_T_72;
  wire [31:0] _GEN_2365 = {{29'd0}, _csrRD_T_74};
  wire [31:0] _csrRD_T_102 = _csrRD_T_100 | _GEN_2365;
  wire [31:0] _csrRD_T_103 = _csrRD_T_102 | _csrRD_T_75;
  wire [31:0] _csrRD_T_104 = _csrRD_T_103 | _csrRD_T_76;
  wire [31:0] csrRD = _csrRD_T_104 | _csrRD_T_77;
  wire [31:0] csrMask = j == 5'h1 ? 32'hffffffff : rj;
  wire [31:0] _crmd_T = rkd & csrMask;
  wire [31:0] _crmd_T_2 = ~csrMask;
  wire [31:0] _GEN_2366 = {{23'd0}, _csrRD_T_1};
  wire [31:0] _crmd_T_3 = _GEN_2366 & _crmd_T_2;
  wire [31:0] _crmd_T_4 = _crmd_T | _crmd_T_3;
  wire  _GEN_182 = _csrRD_T ? _crmd_T_4[4] : crmd_PG;
  wire  _GEN_183 = _csrRD_T ? _crmd_T_4[3] : crmd_DA;
  wire  _GEN_184 = _csrRD_T ? _crmd_T_4[2] : crmd_IE;
  wire [1:0] _GEN_185 = _csrRD_T ? _crmd_T_4[1:0] : crmd_PLV;
  wire [31:0] _GEN_2367 = {{29'd0}, _csrRD_T_3};
  wire [31:0] _prmd_T_3 = _GEN_2367 & _crmd_T_2;
  wire [31:0] _prmd_T_4 = _crmd_T | _prmd_T_3;
  wire  _GEN_186 = _csrRD_T_2 ? _prmd_T_4[2] : csrs_1_PIE;
  wire [1:0] _GEN_187 = _csrRD_T_2 ? _prmd_T_4[1:0] : csrs_1_PPLV;
  wire [31:0] _GEN_2368 = {{31'd0}, csrs_2_FPE};
  wire [31:0] _euen_T_2 = _GEN_2368 & _crmd_T_2;
  wire [31:0] _euen_T_3 = _crmd_T | _euen_T_2;
  wire [31:0] _T_1368 = csrMask & 32'h1bff;
  wire [31:0] _ectl_T = rkd & _T_1368;
  wire [31:0] _ectl_T_1 = ~_T_1368;
  wire [31:0] _GEN_2369 = {{19'd0}, csrs_3_LIE};
  wire [31:0] _ectl_T_2 = _GEN_2369 & _ectl_T_1;
  wire [31:0] _ectl_T_3 = _ectl_T | _ectl_T_2;
  wire [31:0] _era_T_2 = csrs_5_PC & _crmd_T_2;
  wire [31:0] _era_T_3 = _crmd_T | _era_T_2;
  wire [31:0] _GEN_194 = _csrRD_T_8 ? _era_T_3 : csrs_5_PC;
  wire [31:0] _badv_T_2 = badv_VAddr & _crmd_T_2;
  wire [31:0] _badv_T_3 = _crmd_T | _badv_T_2;
  wire [25:0] _eentry_VA_T = rkd[31:6] & csrMask[31:6];
  wire [25:0] _eentry_VA_T_1 = ~csrMask[31:6];
  wire [25:0] _eentry_VA_T_2 = csrs_7_VA & _eentry_VA_T_1;
  wire [25:0] _eentry_VA_T_3 = _eentry_VA_T | _eentry_VA_T_2;
  wire [5:0] _tlbidx_PS_T = rkd[29:24] & csrMask[29:24];
  wire [5:0] _tlbidx_PS_T_1 = ~csrMask[29:24];
  wire [5:0] _tlbidx_PS_T_2 = csrs_8_PS & _tlbidx_PS_T_1;
  wire [5:0] _tlbidx_PS_T_3 = _tlbidx_PS_T | _tlbidx_PS_T_2;
  wire [3:0] _tlbidx_Index_T = rkd[3:0] & csrMask[3:0];
  wire [3:0] _tlbidx_Index_T_1 = ~csrMask[3:0];
  wire [3:0] _tlbidx_Index_T_2 = csrs_8_Index & _tlbidx_Index_T_1;
  wire [3:0] _tlbidx_Index_T_3 = _tlbidx_Index_T | _tlbidx_Index_T_2;
  wire  _GEN_197 = _csrRD_T_12 ? rkd[31] & csrMask[31] | csrs_8_NE & ~csrMask[31] : csrs_8_NE;
  wire [5:0] _GEN_198 = _csrRD_T_12 ? _tlbidx_PS_T_3 : csrs_8_PS;
  wire [3:0] _GEN_199 = _csrRD_T_12 ? _tlbidx_Index_T_3 : csrs_8_Index;
  wire [18:0] _tlbehi_VPPN_T_2 = rkd[31:13] & csrMask[31:13];
  wire [18:0] _tlbehi_VPPN_T_3 = ~csrMask[31:13];
  wire [18:0] _tlbehi_VPPN_T_4 = csrs_9_VPPN & _tlbehi_VPPN_T_3;
  wire [18:0] _tlbehi_VPPN_T_5 = _tlbehi_VPPN_T_2 | _tlbehi_VPPN_T_4;
  wire [18:0] _GEN_200 = _csrRD_T_14 ? _tlbehi_VPPN_T_5 : _GEN_177;
  wire [31:0] _tlbelo0_T_3 = _csrRD_T_17 & _crmd_T_2;
  wire [31:0] _tlbelo0_T_4 = _crmd_T | _tlbelo0_T_3;
  wire [23:0] _tlbelo0_PPN_T = rkd[31:8] & csrMask[31:8];
  wire [23:0] _tlbelo0_PPN_T_1 = ~csrMask[31:8];
  wire [23:0] _tlbelo0_PPN_T_2 = csrs_10_PPN & _tlbelo0_PPN_T_1;
  wire [23:0] _tlbelo0_PPN_T_3 = _tlbelo0_PPN_T | _tlbelo0_PPN_T_2;
  wire [23:0] _GEN_201 = _csrRD_T_16 ? _tlbelo0_PPN_T_3 : csrs_10_PPN;
  wire  _GEN_202 = _csrRD_T_16 ? _tlbelo0_T_4[6] : csrs_10_G;
  wire [1:0] _GEN_203 = _csrRD_T_16 ? _tlbelo0_T_4[5:4] : csrs_10_MAT;
  wire [1:0] _GEN_204 = _csrRD_T_16 ? _tlbelo0_T_4[3:2] : csrs_10_PLV;
  wire  _GEN_205 = _csrRD_T_16 ? _tlbelo0_T_4[1] : csrs_10_D;
  wire  _GEN_206 = _csrRD_T_16 ? _tlbelo0_T_4[0] : csrs_10_V;
  wire [31:0] _tlbelo1_T_3 = _csrRD_T_19 & _crmd_T_2;
  wire [31:0] _tlbelo1_T_4 = _crmd_T | _tlbelo1_T_3;
  wire [23:0] _tlbelo1_PPN_T_2 = csrs_11_PPN & _tlbelo0_PPN_T_1;
  wire [23:0] _tlbelo1_PPN_T_3 = _tlbelo0_PPN_T | _tlbelo1_PPN_T_2;
  wire [23:0] _GEN_207 = _csrRD_T_18 ? _tlbelo1_PPN_T_3 : csrs_11_PPN;
  wire  _GEN_208 = _csrRD_T_18 ? _tlbelo1_T_4[6] : csrs_11_G;
  wire [1:0] _GEN_209 = _csrRD_T_18 ? _tlbelo1_T_4[5:4] : csrs_11_MAT;
  wire [1:0] _GEN_210 = _csrRD_T_18 ? _tlbelo1_T_4[3:2] : csrs_11_PLV;
  wire  _GEN_211 = _csrRD_T_18 ? _tlbelo1_T_4[1] : csrs_11_D;
  wire  _GEN_212 = _csrRD_T_18 ? _tlbelo1_T_4[0] : csrs_11_V;
  wire [9:0] _asid_ASID_T = rkd[9:0] & csrMask[9:0];
  wire [9:0] _asid_ASID_T_1 = ~csrMask[9:0];
  wire [9:0] _asid_ASID_T_2 = asid_ASID & _asid_ASID_T_1;
  wire [9:0] _asid_ASID_T_3 = _asid_ASID_T | _asid_ASID_T_2;
  wire [9:0] _GEN_213 = _csrRD_T_20 ? _asid_ASID_T_3 : asid_ASID;
  wire [19:0] _pgdl_Base_T = rkd[31:12] & csrMask[31:12];
  wire [19:0] _pgdl_Base_T_1 = ~csrMask[31:12];
  wire [19:0] _pgdl_Base_T_2 = csrs_13_Base & _pgdl_Base_T_1;
  wire [19:0] _pgdl_Base_T_3 = _pgdl_Base_T | _pgdl_Base_T_2;
  wire [19:0] _pgdh_Base_T_2 = csrs_14_Base & _pgdl_Base_T_1;
  wire [19:0] _pgdh_Base_T_3 = _pgdl_Base_T | _pgdh_Base_T_2;
  wire [31:0] _save0_T_2 = csrs_17_Data & _crmd_T_2;
  wire [31:0] _save0_T_3 = _crmd_T | _save0_T_2;
  wire [31:0] _save1_T_2 = csrs_18_Data & _crmd_T_2;
  wire [31:0] _save1_T_3 = _crmd_T | _save1_T_2;
  wire [31:0] _save2_T_2 = csrs_19_Data & _crmd_T_2;
  wire [31:0] _save2_T_3 = _crmd_T | _save2_T_2;
  wire [31:0] _save3_T_2 = csrs_20_Data & _crmd_T_2;
  wire [31:0] _save3_T_3 = _crmd_T | _save3_T_2;
  wire [31:0] _tid_T_2 = csrs_21_TID & _crmd_T_2;
  wire [31:0] _tid_T_3 = _crmd_T | _tid_T_2;
  wire [31:0] _next_T_3 = _csrRD_T_38 & _crmd_T_2;
  wire [31:0] _next_T_4 = _crmd_T | _next_T_3;
  wire  next_En = _next_T_4[0];
  wire  next_Periodic = _next_T_4[1];
  wire [29:0] next_InitVal = _next_T_4[31:2];
  wire [31:0] _tval_TimeVal_T_3 = {next_InitVal,2'h0};
  wire  _GEN_221 = next_InitVal == 30'h0 | _GEN_5;
  wire  _GEN_223 = next_En ? _GEN_221 : _GEN_5;
  wire  _GEN_228 = _csrRD_T_37 ? _GEN_223 : _GEN_5;
  wire  _T_1415 = rkd[0] & csrMask[0];
  wire  _GEN_231 = csrMask[2] ? rkd[2] : csrs_25_KLO;
  wire  _GEN_232 = csrMask[1] & rkd[1] ? 1'h0 : _GEN_179;
  wire  _GEN_234 = _csrRD_T_41 ? _GEN_232 : _GEN_179;
  wire [25:0] _tlbrentry_PA_T_2 = csrs_26_PA & _eentry_VA_T_1;
  wire [25:0] _tlbrentry_PA_T_3 = _eentry_VA_T | _tlbrentry_PA_T_2;
  wire [1:0] _dmw0_MAT_T = rkd[5:4] & csrMask[5:4];
  wire [1:0] _dmw0_MAT_T_1 = ~csrMask[5:4];
  wire [1:0] _dmw0_MAT_T_2 = csrs_27_MAT & _dmw0_MAT_T_1;
  wire [1:0] _dmw0_MAT_T_3 = _dmw0_MAT_T | _dmw0_MAT_T_2;
  wire [2:0] _dmw0_PSEG_T = rkd[27:25] & csrMask[27:25];
  wire [2:0] _dmw0_PSEG_T_1 = ~csrMask[27:25];
  wire [2:0] _dmw0_PSEG_T_2 = csrs_27_PSEG & _dmw0_PSEG_T_1;
  wire [2:0] _dmw0_PSEG_T_3 = _dmw0_PSEG_T | _dmw0_PSEG_T_2;
  wire [2:0] _dmw0_VSEG_T = rkd[31:29] & csrMask[31:29];
  wire [2:0] _dmw0_VSEG_T_1 = ~csrMask[31:29];
  wire [2:0] _dmw0_VSEG_T_2 = csrs_27_VSEG & _dmw0_VSEG_T_1;
  wire [2:0] _dmw0_VSEG_T_3 = _dmw0_VSEG_T | _dmw0_VSEG_T_2;
  wire [1:0] _dmw1_MAT_T_2 = csrs_28_MAT & _dmw0_MAT_T_1;
  wire [1:0] _dmw1_MAT_T_3 = _dmw0_MAT_T | _dmw1_MAT_T_2;
  wire [2:0] _dmw1_PSEG_T_2 = csrs_28_PSEG & _dmw0_PSEG_T_1;
  wire [2:0] _dmw1_PSEG_T_3 = _dmw0_PSEG_T | _dmw1_PSEG_T_2;
  wire [2:0] _dmw1_VSEG_T_2 = csrs_28_VSEG & _dmw0_VSEG_T_1;
  wire [2:0] _dmw1_VSEG_T_3 = _dmw0_VSEG_T | _dmw1_VSEG_T_2;
  wire  _GEN_248 = ID_OK & c0_4 & |csrMask ? _GEN_182 : crmd_PG;
  wire  _GEN_249 = ID_OK & c0_4 & |csrMask ? _GEN_183 : crmd_DA;
  wire  _GEN_250 = ID_OK & c0_4 & |csrMask ? _GEN_184 : crmd_IE;
  wire [1:0] _GEN_251 = ID_OK & c0_4 & |csrMask ? _GEN_185 : crmd_PLV;
  wire  _GEN_252 = ID_OK & c0_4 & |csrMask ? _GEN_186 : csrs_1_PIE;
  wire [1:0] _GEN_253 = ID_OK & c0_4 & |csrMask ? _GEN_187 : csrs_1_PPLV;
  wire [31:0] _GEN_258 = ID_OK & c0_4 & |csrMask ? _GEN_194 : csrs_5_PC;
  wire  _GEN_261 = ID_OK & c0_4 & |csrMask ? _GEN_197 : csrs_8_NE;
  wire [5:0] _GEN_262 = ID_OK & c0_4 & |csrMask ? _GEN_198 : csrs_8_PS;
  wire [3:0] _GEN_263 = ID_OK & c0_4 & |csrMask ? _GEN_199 : csrs_8_Index;
  wire [18:0] _GEN_264 = ID_OK & c0_4 & |csrMask ? _GEN_200 : _GEN_177;
  wire [23:0] _GEN_265 = ID_OK & c0_4 & |csrMask ? _GEN_201 : csrs_10_PPN;
  wire  _GEN_266 = ID_OK & c0_4 & |csrMask ? _GEN_202 : csrs_10_G;
  wire [1:0] _GEN_267 = ID_OK & c0_4 & |csrMask ? _GEN_203 : csrs_10_MAT;
  wire [1:0] _GEN_268 = ID_OK & c0_4 & |csrMask ? _GEN_204 : csrs_10_PLV;
  wire  _GEN_269 = ID_OK & c0_4 & |csrMask ? _GEN_205 : csrs_10_D;
  wire  _GEN_270 = ID_OK & c0_4 & |csrMask ? _GEN_206 : csrs_10_V;
  wire [23:0] _GEN_271 = ID_OK & c0_4 & |csrMask ? _GEN_207 : csrs_11_PPN;
  wire  _GEN_272 = ID_OK & c0_4 & |csrMask ? _GEN_208 : csrs_11_G;
  wire [1:0] _GEN_273 = ID_OK & c0_4 & |csrMask ? _GEN_209 : csrs_11_MAT;
  wire [1:0] _GEN_274 = ID_OK & c0_4 & |csrMask ? _GEN_210 : csrs_11_PLV;
  wire  _GEN_275 = ID_OK & c0_4 & |csrMask ? _GEN_211 : csrs_11_D;
  wire  _GEN_276 = ID_OK & c0_4 & |csrMask ? _GEN_212 : csrs_11_V;
  wire [9:0] _GEN_277 = ID_OK & c0_4 & |csrMask ? _GEN_213 : asid_ASID;
  wire  _GEN_291 = ID_OK & c0_4 & |csrMask ? _GEN_234 : _GEN_179;
  wire [3:0] _tlbidx_Index_T_5 = tlbHit_1_1 ? 4'h1 : 4'h0;
  wire [3:0] _tlbidx_Index_T_6 = tlbHit_2_1 ? 4'h2 : 4'h0;
  wire [3:0] _tlbidx_Index_T_7 = tlbHit_3_1 ? 4'h3 : 4'h0;
  wire [3:0] _tlbidx_Index_T_8 = tlbHit_4_1 ? 4'h4 : 4'h0;
  wire [3:0] _tlbidx_Index_T_9 = tlbHit_5_1 ? 4'h5 : 4'h0;
  wire [3:0] _tlbidx_Index_T_10 = tlbHit_6_1 ? 4'h6 : 4'h0;
  wire [3:0] _tlbidx_Index_T_11 = tlbHit_7_1 ? 4'h7 : 4'h0;
  wire [3:0] _tlbidx_Index_T_12 = tlbHit_8_1 ? 4'h8 : 4'h0;
  wire [3:0] _tlbidx_Index_T_13 = tlbHit_9_1 ? 4'h9 : 4'h0;
  wire [3:0] _tlbidx_Index_T_14 = tlbHit_10_1 ? 4'ha : 4'h0;
  wire [3:0] _tlbidx_Index_T_15 = tlbHit_11_1 ? 4'hb : 4'h0;
  wire [3:0] _tlbidx_Index_T_16 = tlbHit_12_1 ? 4'hc : 4'h0;
  wire [3:0] _tlbidx_Index_T_17 = tlbHit_13_1 ? 4'hd : 4'h0;
  wire [3:0] _tlbidx_Index_T_18 = tlbHit_14_1 ? 4'he : 4'h0;
  wire [3:0] _tlbidx_Index_T_19 = tlbHit_15_1 ? 4'hf : 4'h0;
  wire [3:0] _tlbidx_Index_T_21 = _tlbidx_Index_T_5 | _tlbidx_Index_T_6;
  wire [3:0] _tlbidx_Index_T_22 = _tlbidx_Index_T_21 | _tlbidx_Index_T_7;
  wire [3:0] _tlbidx_Index_T_23 = _tlbidx_Index_T_22 | _tlbidx_Index_T_8;
  wire [3:0] _tlbidx_Index_T_24 = _tlbidx_Index_T_23 | _tlbidx_Index_T_9;
  wire [3:0] _tlbidx_Index_T_25 = _tlbidx_Index_T_24 | _tlbidx_Index_T_10;
  wire [3:0] _tlbidx_Index_T_26 = _tlbidx_Index_T_25 | _tlbidx_Index_T_11;
  wire [3:0] _tlbidx_Index_T_27 = _tlbidx_Index_T_26 | _tlbidx_Index_T_12;
  wire [3:0] _tlbidx_Index_T_28 = _tlbidx_Index_T_27 | _tlbidx_Index_T_13;
  wire [3:0] _tlbidx_Index_T_29 = _tlbidx_Index_T_28 | _tlbidx_Index_T_14;
  wire [3:0] _tlbidx_Index_T_30 = _tlbidx_Index_T_29 | _tlbidx_Index_T_15;
  wire [3:0] _tlbidx_Index_T_31 = _tlbidx_Index_T_30 | _tlbidx_Index_T_16;
  wire [3:0] _tlbidx_Index_T_32 = _tlbidx_Index_T_31 | _tlbidx_Index_T_17;
  wire [3:0] _tlbidx_Index_T_33 = _tlbidx_Index_T_32 | _tlbidx_Index_T_18;
  wire [3:0] _tlbidx_Index_T_34 = _tlbidx_Index_T_33 | _tlbidx_Index_T_19;
  wire  _GEN_306 = 4'h1 == csrs_8_Index ? tlb_1_E : tlb_0_E;
  wire  _GEN_307 = 4'h2 == csrs_8_Index ? tlb_2_E : _GEN_306;
  wire  _GEN_308 = 4'h3 == csrs_8_Index ? tlb_3_E : _GEN_307;
  wire  _GEN_309 = 4'h4 == csrs_8_Index ? tlb_4_E : _GEN_308;
  wire  _GEN_310 = 4'h5 == csrs_8_Index ? tlb_5_E : _GEN_309;
  wire  _GEN_311 = 4'h6 == csrs_8_Index ? tlb_6_E : _GEN_310;
  wire  _GEN_312 = 4'h7 == csrs_8_Index ? tlb_7_E : _GEN_311;
  wire  _GEN_313 = 4'h8 == csrs_8_Index ? tlb_8_E : _GEN_312;
  wire  _GEN_314 = 4'h9 == csrs_8_Index ? tlb_9_E : _GEN_313;
  wire  _GEN_315 = 4'ha == csrs_8_Index ? tlb_10_E : _GEN_314;
  wire  _GEN_316 = 4'hb == csrs_8_Index ? tlb_11_E : _GEN_315;
  wire  _GEN_317 = 4'hc == csrs_8_Index ? tlb_12_E : _GEN_316;
  wire  _GEN_318 = 4'hd == csrs_8_Index ? tlb_13_E : _GEN_317;
  wire  _GEN_319 = 4'he == csrs_8_Index ? tlb_14_E : _GEN_318;
  wire  _GEN_320 = 4'hf == csrs_8_Index ? tlb_15_E : _GEN_319;
  wire [5:0] _GEN_322 = 4'h1 == csrs_8_Index ? tlb_1_PS : tlb_0_PS;
  wire [5:0] _GEN_323 = 4'h2 == csrs_8_Index ? tlb_2_PS : _GEN_322;
  wire [5:0] _GEN_324 = 4'h3 == csrs_8_Index ? tlb_3_PS : _GEN_323;
  wire [5:0] _GEN_325 = 4'h4 == csrs_8_Index ? tlb_4_PS : _GEN_324;
  wire [5:0] _GEN_326 = 4'h5 == csrs_8_Index ? tlb_5_PS : _GEN_325;
  wire [5:0] _GEN_327 = 4'h6 == csrs_8_Index ? tlb_6_PS : _GEN_326;
  wire [5:0] _GEN_328 = 4'h7 == csrs_8_Index ? tlb_7_PS : _GEN_327;
  wire [5:0] _GEN_329 = 4'h8 == csrs_8_Index ? tlb_8_PS : _GEN_328;
  wire [5:0] _GEN_330 = 4'h9 == csrs_8_Index ? tlb_9_PS : _GEN_329;
  wire [5:0] _GEN_331 = 4'ha == csrs_8_Index ? tlb_10_PS : _GEN_330;
  wire [5:0] _GEN_332 = 4'hb == csrs_8_Index ? tlb_11_PS : _GEN_331;
  wire [5:0] _GEN_333 = 4'hc == csrs_8_Index ? tlb_12_PS : _GEN_332;
  wire [5:0] _GEN_334 = 4'hd == csrs_8_Index ? tlb_13_PS : _GEN_333;
  wire [5:0] _GEN_335 = 4'he == csrs_8_Index ? tlb_14_PS : _GEN_334;
  wire [5:0] _GEN_336 = 4'hf == csrs_8_Index ? tlb_15_PS : _GEN_335;
  wire [18:0] _GEN_338 = 4'h1 == csrs_8_Index ? tlb_1_VPPN : tlb_0_VPPN;
  wire [18:0] _GEN_339 = 4'h2 == csrs_8_Index ? tlb_2_VPPN : _GEN_338;
  wire [18:0] _GEN_340 = 4'h3 == csrs_8_Index ? tlb_3_VPPN : _GEN_339;
  wire [18:0] _GEN_341 = 4'h4 == csrs_8_Index ? tlb_4_VPPN : _GEN_340;
  wire [18:0] _GEN_342 = 4'h5 == csrs_8_Index ? tlb_5_VPPN : _GEN_341;
  wire [18:0] _GEN_343 = 4'h6 == csrs_8_Index ? tlb_6_VPPN : _GEN_342;
  wire [18:0] _GEN_344 = 4'h7 == csrs_8_Index ? tlb_7_VPPN : _GEN_343;
  wire [18:0] _GEN_345 = 4'h8 == csrs_8_Index ? tlb_8_VPPN : _GEN_344;
  wire [18:0] _GEN_346 = 4'h9 == csrs_8_Index ? tlb_9_VPPN : _GEN_345;
  wire [18:0] _GEN_347 = 4'ha == csrs_8_Index ? tlb_10_VPPN : _GEN_346;
  wire [18:0] _GEN_348 = 4'hb == csrs_8_Index ? tlb_11_VPPN : _GEN_347;
  wire [18:0] _GEN_349 = 4'hc == csrs_8_Index ? tlb_12_VPPN : _GEN_348;
  wire [18:0] _GEN_350 = 4'hd == csrs_8_Index ? tlb_13_VPPN : _GEN_349;
  wire [18:0] _GEN_351 = 4'he == csrs_8_Index ? tlb_14_VPPN : _GEN_350;
  wire [18:0] _GEN_352 = 4'hf == csrs_8_Index ? tlb_15_VPPN : _GEN_351;
  wire [19:0] _GEN_354 = 4'h1 == csrs_8_Index ? tlb_1_P0_PPN : tlb_0_P0_PPN;
  wire [19:0] _GEN_355 = 4'h2 == csrs_8_Index ? tlb_2_P0_PPN : _GEN_354;
  wire [19:0] _GEN_356 = 4'h3 == csrs_8_Index ? tlb_3_P0_PPN : _GEN_355;
  wire [19:0] _GEN_357 = 4'h4 == csrs_8_Index ? tlb_4_P0_PPN : _GEN_356;
  wire [19:0] _GEN_358 = 4'h5 == csrs_8_Index ? tlb_5_P0_PPN : _GEN_357;
  wire [19:0] _GEN_359 = 4'h6 == csrs_8_Index ? tlb_6_P0_PPN : _GEN_358;
  wire [19:0] _GEN_360 = 4'h7 == csrs_8_Index ? tlb_7_P0_PPN : _GEN_359;
  wire [19:0] _GEN_361 = 4'h8 == csrs_8_Index ? tlb_8_P0_PPN : _GEN_360;
  wire [19:0] _GEN_362 = 4'h9 == csrs_8_Index ? tlb_9_P0_PPN : _GEN_361;
  wire [19:0] _GEN_363 = 4'ha == csrs_8_Index ? tlb_10_P0_PPN : _GEN_362;
  wire [19:0] _GEN_364 = 4'hb == csrs_8_Index ? tlb_11_P0_PPN : _GEN_363;
  wire [19:0] _GEN_365 = 4'hc == csrs_8_Index ? tlb_12_P0_PPN : _GEN_364;
  wire [19:0] _GEN_366 = 4'hd == csrs_8_Index ? tlb_13_P0_PPN : _GEN_365;
  wire [19:0] _GEN_367 = 4'he == csrs_8_Index ? tlb_14_P0_PPN : _GEN_366;
  wire [19:0] _GEN_368 = 4'hf == csrs_8_Index ? tlb_15_P0_PPN : _GEN_367;
  wire  _GEN_370 = 4'h1 == csrs_8_Index ? tlb_1_G : tlb_0_G;
  wire  _GEN_371 = 4'h2 == csrs_8_Index ? tlb_2_G : _GEN_370;
  wire  _GEN_372 = 4'h3 == csrs_8_Index ? tlb_3_G : _GEN_371;
  wire  _GEN_373 = 4'h4 == csrs_8_Index ? tlb_4_G : _GEN_372;
  wire  _GEN_374 = 4'h5 == csrs_8_Index ? tlb_5_G : _GEN_373;
  wire  _GEN_375 = 4'h6 == csrs_8_Index ? tlb_6_G : _GEN_374;
  wire  _GEN_376 = 4'h7 == csrs_8_Index ? tlb_7_G : _GEN_375;
  wire  _GEN_377 = 4'h8 == csrs_8_Index ? tlb_8_G : _GEN_376;
  wire  _GEN_378 = 4'h9 == csrs_8_Index ? tlb_9_G : _GEN_377;
  wire  _GEN_379 = 4'ha == csrs_8_Index ? tlb_10_G : _GEN_378;
  wire  _GEN_380 = 4'hb == csrs_8_Index ? tlb_11_G : _GEN_379;
  wire  _GEN_381 = 4'hc == csrs_8_Index ? tlb_12_G : _GEN_380;
  wire  _GEN_382 = 4'hd == csrs_8_Index ? tlb_13_G : _GEN_381;
  wire  _GEN_383 = 4'he == csrs_8_Index ? tlb_14_G : _GEN_382;
  wire  _GEN_384 = 4'hf == csrs_8_Index ? tlb_15_G : _GEN_383;
  wire [1:0] _GEN_386 = 4'h1 == csrs_8_Index ? tlb_1_P0_MAT : tlb_0_P0_MAT;
  wire [1:0] _GEN_387 = 4'h2 == csrs_8_Index ? tlb_2_P0_MAT : _GEN_386;
  wire [1:0] _GEN_388 = 4'h3 == csrs_8_Index ? tlb_3_P0_MAT : _GEN_387;
  wire [1:0] _GEN_389 = 4'h4 == csrs_8_Index ? tlb_4_P0_MAT : _GEN_388;
  wire [1:0] _GEN_390 = 4'h5 == csrs_8_Index ? tlb_5_P0_MAT : _GEN_389;
  wire [1:0] _GEN_391 = 4'h6 == csrs_8_Index ? tlb_6_P0_MAT : _GEN_390;
  wire [1:0] _GEN_392 = 4'h7 == csrs_8_Index ? tlb_7_P0_MAT : _GEN_391;
  wire [1:0] _GEN_393 = 4'h8 == csrs_8_Index ? tlb_8_P0_MAT : _GEN_392;
  wire [1:0] _GEN_394 = 4'h9 == csrs_8_Index ? tlb_9_P0_MAT : _GEN_393;
  wire [1:0] _GEN_395 = 4'ha == csrs_8_Index ? tlb_10_P0_MAT : _GEN_394;
  wire [1:0] _GEN_396 = 4'hb == csrs_8_Index ? tlb_11_P0_MAT : _GEN_395;
  wire [1:0] _GEN_397 = 4'hc == csrs_8_Index ? tlb_12_P0_MAT : _GEN_396;
  wire [1:0] _GEN_398 = 4'hd == csrs_8_Index ? tlb_13_P0_MAT : _GEN_397;
  wire [1:0] _GEN_399 = 4'he == csrs_8_Index ? tlb_14_P0_MAT : _GEN_398;
  wire [1:0] _GEN_400 = 4'hf == csrs_8_Index ? tlb_15_P0_MAT : _GEN_399;
  wire [1:0] _GEN_402 = 4'h1 == csrs_8_Index ? tlb_1_P0_PLV : tlb_0_P0_PLV;
  wire [1:0] _GEN_403 = 4'h2 == csrs_8_Index ? tlb_2_P0_PLV : _GEN_402;
  wire [1:0] _GEN_404 = 4'h3 == csrs_8_Index ? tlb_3_P0_PLV : _GEN_403;
  wire [1:0] _GEN_405 = 4'h4 == csrs_8_Index ? tlb_4_P0_PLV : _GEN_404;
  wire [1:0] _GEN_406 = 4'h5 == csrs_8_Index ? tlb_5_P0_PLV : _GEN_405;
  wire [1:0] _GEN_407 = 4'h6 == csrs_8_Index ? tlb_6_P0_PLV : _GEN_406;
  wire [1:0] _GEN_408 = 4'h7 == csrs_8_Index ? tlb_7_P0_PLV : _GEN_407;
  wire [1:0] _GEN_409 = 4'h8 == csrs_8_Index ? tlb_8_P0_PLV : _GEN_408;
  wire [1:0] _GEN_410 = 4'h9 == csrs_8_Index ? tlb_9_P0_PLV : _GEN_409;
  wire [1:0] _GEN_411 = 4'ha == csrs_8_Index ? tlb_10_P0_PLV : _GEN_410;
  wire [1:0] _GEN_412 = 4'hb == csrs_8_Index ? tlb_11_P0_PLV : _GEN_411;
  wire [1:0] _GEN_413 = 4'hc == csrs_8_Index ? tlb_12_P0_PLV : _GEN_412;
  wire [1:0] _GEN_414 = 4'hd == csrs_8_Index ? tlb_13_P0_PLV : _GEN_413;
  wire [1:0] _GEN_415 = 4'he == csrs_8_Index ? tlb_14_P0_PLV : _GEN_414;
  wire [1:0] _GEN_416 = 4'hf == csrs_8_Index ? tlb_15_P0_PLV : _GEN_415;
  wire  _GEN_418 = 4'h1 == csrs_8_Index ? tlb_1_P0_D : tlb_0_P0_D;
  wire  _GEN_419 = 4'h2 == csrs_8_Index ? tlb_2_P0_D : _GEN_418;
  wire  _GEN_420 = 4'h3 == csrs_8_Index ? tlb_3_P0_D : _GEN_419;
  wire  _GEN_421 = 4'h4 == csrs_8_Index ? tlb_4_P0_D : _GEN_420;
  wire  _GEN_422 = 4'h5 == csrs_8_Index ? tlb_5_P0_D : _GEN_421;
  wire  _GEN_423 = 4'h6 == csrs_8_Index ? tlb_6_P0_D : _GEN_422;
  wire  _GEN_424 = 4'h7 == csrs_8_Index ? tlb_7_P0_D : _GEN_423;
  wire  _GEN_425 = 4'h8 == csrs_8_Index ? tlb_8_P0_D : _GEN_424;
  wire  _GEN_426 = 4'h9 == csrs_8_Index ? tlb_9_P0_D : _GEN_425;
  wire  _GEN_427 = 4'ha == csrs_8_Index ? tlb_10_P0_D : _GEN_426;
  wire  _GEN_428 = 4'hb == csrs_8_Index ? tlb_11_P0_D : _GEN_427;
  wire  _GEN_429 = 4'hc == csrs_8_Index ? tlb_12_P0_D : _GEN_428;
  wire  _GEN_430 = 4'hd == csrs_8_Index ? tlb_13_P0_D : _GEN_429;
  wire  _GEN_431 = 4'he == csrs_8_Index ? tlb_14_P0_D : _GEN_430;
  wire  _GEN_432 = 4'hf == csrs_8_Index ? tlb_15_P0_D : _GEN_431;
  wire  _GEN_434 = 4'h1 == csrs_8_Index ? tlb_1_P0_V : tlb_0_P0_V;
  wire  _GEN_435 = 4'h2 == csrs_8_Index ? tlb_2_P0_V : _GEN_434;
  wire  _GEN_436 = 4'h3 == csrs_8_Index ? tlb_3_P0_V : _GEN_435;
  wire  _GEN_437 = 4'h4 == csrs_8_Index ? tlb_4_P0_V : _GEN_436;
  wire  _GEN_438 = 4'h5 == csrs_8_Index ? tlb_5_P0_V : _GEN_437;
  wire  _GEN_439 = 4'h6 == csrs_8_Index ? tlb_6_P0_V : _GEN_438;
  wire  _GEN_440 = 4'h7 == csrs_8_Index ? tlb_7_P0_V : _GEN_439;
  wire  _GEN_441 = 4'h8 == csrs_8_Index ? tlb_8_P0_V : _GEN_440;
  wire  _GEN_442 = 4'h9 == csrs_8_Index ? tlb_9_P0_V : _GEN_441;
  wire  _GEN_443 = 4'ha == csrs_8_Index ? tlb_10_P0_V : _GEN_442;
  wire  _GEN_444 = 4'hb == csrs_8_Index ? tlb_11_P0_V : _GEN_443;
  wire  _GEN_445 = 4'hc == csrs_8_Index ? tlb_12_P0_V : _GEN_444;
  wire  _GEN_446 = 4'hd == csrs_8_Index ? tlb_13_P0_V : _GEN_445;
  wire  _GEN_447 = 4'he == csrs_8_Index ? tlb_14_P0_V : _GEN_446;
  wire  _GEN_448 = 4'hf == csrs_8_Index ? tlb_15_P0_V : _GEN_447;
  wire [19:0] _GEN_450 = 4'h1 == csrs_8_Index ? tlb_1_P1_PPN : tlb_0_P1_PPN;
  wire [19:0] _GEN_451 = 4'h2 == csrs_8_Index ? tlb_2_P1_PPN : _GEN_450;
  wire [19:0] _GEN_452 = 4'h3 == csrs_8_Index ? tlb_3_P1_PPN : _GEN_451;
  wire [19:0] _GEN_453 = 4'h4 == csrs_8_Index ? tlb_4_P1_PPN : _GEN_452;
  wire [19:0] _GEN_454 = 4'h5 == csrs_8_Index ? tlb_5_P1_PPN : _GEN_453;
  wire [19:0] _GEN_455 = 4'h6 == csrs_8_Index ? tlb_6_P1_PPN : _GEN_454;
  wire [19:0] _GEN_456 = 4'h7 == csrs_8_Index ? tlb_7_P1_PPN : _GEN_455;
  wire [19:0] _GEN_457 = 4'h8 == csrs_8_Index ? tlb_8_P1_PPN : _GEN_456;
  wire [19:0] _GEN_458 = 4'h9 == csrs_8_Index ? tlb_9_P1_PPN : _GEN_457;
  wire [19:0] _GEN_459 = 4'ha == csrs_8_Index ? tlb_10_P1_PPN : _GEN_458;
  wire [19:0] _GEN_460 = 4'hb == csrs_8_Index ? tlb_11_P1_PPN : _GEN_459;
  wire [19:0] _GEN_461 = 4'hc == csrs_8_Index ? tlb_12_P1_PPN : _GEN_460;
  wire [19:0] _GEN_462 = 4'hd == csrs_8_Index ? tlb_13_P1_PPN : _GEN_461;
  wire [19:0] _GEN_463 = 4'he == csrs_8_Index ? tlb_14_P1_PPN : _GEN_462;
  wire [19:0] _GEN_464 = 4'hf == csrs_8_Index ? tlb_15_P1_PPN : _GEN_463;
  wire [1:0] _GEN_466 = 4'h1 == csrs_8_Index ? tlb_1_P1_MAT : tlb_0_P1_MAT;
  wire [1:0] _GEN_467 = 4'h2 == csrs_8_Index ? tlb_2_P1_MAT : _GEN_466;
  wire [1:0] _GEN_468 = 4'h3 == csrs_8_Index ? tlb_3_P1_MAT : _GEN_467;
  wire [1:0] _GEN_469 = 4'h4 == csrs_8_Index ? tlb_4_P1_MAT : _GEN_468;
  wire [1:0] _GEN_470 = 4'h5 == csrs_8_Index ? tlb_5_P1_MAT : _GEN_469;
  wire [1:0] _GEN_471 = 4'h6 == csrs_8_Index ? tlb_6_P1_MAT : _GEN_470;
  wire [1:0] _GEN_472 = 4'h7 == csrs_8_Index ? tlb_7_P1_MAT : _GEN_471;
  wire [1:0] _GEN_473 = 4'h8 == csrs_8_Index ? tlb_8_P1_MAT : _GEN_472;
  wire [1:0] _GEN_474 = 4'h9 == csrs_8_Index ? tlb_9_P1_MAT : _GEN_473;
  wire [1:0] _GEN_475 = 4'ha == csrs_8_Index ? tlb_10_P1_MAT : _GEN_474;
  wire [1:0] _GEN_476 = 4'hb == csrs_8_Index ? tlb_11_P1_MAT : _GEN_475;
  wire [1:0] _GEN_477 = 4'hc == csrs_8_Index ? tlb_12_P1_MAT : _GEN_476;
  wire [1:0] _GEN_478 = 4'hd == csrs_8_Index ? tlb_13_P1_MAT : _GEN_477;
  wire [1:0] _GEN_479 = 4'he == csrs_8_Index ? tlb_14_P1_MAT : _GEN_478;
  wire [1:0] _GEN_480 = 4'hf == csrs_8_Index ? tlb_15_P1_MAT : _GEN_479;
  wire [1:0] _GEN_482 = 4'h1 == csrs_8_Index ? tlb_1_P1_PLV : tlb_0_P1_PLV;
  wire [1:0] _GEN_483 = 4'h2 == csrs_8_Index ? tlb_2_P1_PLV : _GEN_482;
  wire [1:0] _GEN_484 = 4'h3 == csrs_8_Index ? tlb_3_P1_PLV : _GEN_483;
  wire [1:0] _GEN_485 = 4'h4 == csrs_8_Index ? tlb_4_P1_PLV : _GEN_484;
  wire [1:0] _GEN_486 = 4'h5 == csrs_8_Index ? tlb_5_P1_PLV : _GEN_485;
  wire [1:0] _GEN_487 = 4'h6 == csrs_8_Index ? tlb_6_P1_PLV : _GEN_486;
  wire [1:0] _GEN_488 = 4'h7 == csrs_8_Index ? tlb_7_P1_PLV : _GEN_487;
  wire [1:0] _GEN_489 = 4'h8 == csrs_8_Index ? tlb_8_P1_PLV : _GEN_488;
  wire [1:0] _GEN_490 = 4'h9 == csrs_8_Index ? tlb_9_P1_PLV : _GEN_489;
  wire [1:0] _GEN_491 = 4'ha == csrs_8_Index ? tlb_10_P1_PLV : _GEN_490;
  wire [1:0] _GEN_492 = 4'hb == csrs_8_Index ? tlb_11_P1_PLV : _GEN_491;
  wire [1:0] _GEN_493 = 4'hc == csrs_8_Index ? tlb_12_P1_PLV : _GEN_492;
  wire [1:0] _GEN_494 = 4'hd == csrs_8_Index ? tlb_13_P1_PLV : _GEN_493;
  wire [1:0] _GEN_495 = 4'he == csrs_8_Index ? tlb_14_P1_PLV : _GEN_494;
  wire [1:0] _GEN_496 = 4'hf == csrs_8_Index ? tlb_15_P1_PLV : _GEN_495;
  wire  _GEN_498 = 4'h1 == csrs_8_Index ? tlb_1_P1_D : tlb_0_P1_D;
  wire  _GEN_499 = 4'h2 == csrs_8_Index ? tlb_2_P1_D : _GEN_498;
  wire  _GEN_500 = 4'h3 == csrs_8_Index ? tlb_3_P1_D : _GEN_499;
  wire  _GEN_501 = 4'h4 == csrs_8_Index ? tlb_4_P1_D : _GEN_500;
  wire  _GEN_502 = 4'h5 == csrs_8_Index ? tlb_5_P1_D : _GEN_501;
  wire  _GEN_503 = 4'h6 == csrs_8_Index ? tlb_6_P1_D : _GEN_502;
  wire  _GEN_504 = 4'h7 == csrs_8_Index ? tlb_7_P1_D : _GEN_503;
  wire  _GEN_505 = 4'h8 == csrs_8_Index ? tlb_8_P1_D : _GEN_504;
  wire  _GEN_506 = 4'h9 == csrs_8_Index ? tlb_9_P1_D : _GEN_505;
  wire  _GEN_507 = 4'ha == csrs_8_Index ? tlb_10_P1_D : _GEN_506;
  wire  _GEN_508 = 4'hb == csrs_8_Index ? tlb_11_P1_D : _GEN_507;
  wire  _GEN_509 = 4'hc == csrs_8_Index ? tlb_12_P1_D : _GEN_508;
  wire  _GEN_510 = 4'hd == csrs_8_Index ? tlb_13_P1_D : _GEN_509;
  wire  _GEN_511 = 4'he == csrs_8_Index ? tlb_14_P1_D : _GEN_510;
  wire  _GEN_512 = 4'hf == csrs_8_Index ? tlb_15_P1_D : _GEN_511;
  wire  _GEN_514 = 4'h1 == csrs_8_Index ? tlb_1_P1_V : tlb_0_P1_V;
  wire  _GEN_515 = 4'h2 == csrs_8_Index ? tlb_2_P1_V : _GEN_514;
  wire  _GEN_516 = 4'h3 == csrs_8_Index ? tlb_3_P1_V : _GEN_515;
  wire  _GEN_517 = 4'h4 == csrs_8_Index ? tlb_4_P1_V : _GEN_516;
  wire  _GEN_518 = 4'h5 == csrs_8_Index ? tlb_5_P1_V : _GEN_517;
  wire  _GEN_519 = 4'h6 == csrs_8_Index ? tlb_6_P1_V : _GEN_518;
  wire  _GEN_520 = 4'h7 == csrs_8_Index ? tlb_7_P1_V : _GEN_519;
  wire  _GEN_521 = 4'h8 == csrs_8_Index ? tlb_8_P1_V : _GEN_520;
  wire  _GEN_522 = 4'h9 == csrs_8_Index ? tlb_9_P1_V : _GEN_521;
  wire  _GEN_523 = 4'ha == csrs_8_Index ? tlb_10_P1_V : _GEN_522;
  wire  _GEN_524 = 4'hb == csrs_8_Index ? tlb_11_P1_V : _GEN_523;
  wire  _GEN_525 = 4'hc == csrs_8_Index ? tlb_12_P1_V : _GEN_524;
  wire  _GEN_526 = 4'hd == csrs_8_Index ? tlb_13_P1_V : _GEN_525;
  wire  _GEN_527 = 4'he == csrs_8_Index ? tlb_14_P1_V : _GEN_526;
  wire  _GEN_528 = 4'hf == csrs_8_Index ? tlb_15_P1_V : _GEN_527;
  wire [9:0] _GEN_530 = 4'h1 == csrs_8_Index ? tlb_1_ASID : tlb_0_ASID;
  wire [9:0] _GEN_531 = 4'h2 == csrs_8_Index ? tlb_2_ASID : _GEN_530;
  wire [9:0] _GEN_532 = 4'h3 == csrs_8_Index ? tlb_3_ASID : _GEN_531;
  wire [9:0] _GEN_533 = 4'h4 == csrs_8_Index ? tlb_4_ASID : _GEN_532;
  wire [9:0] _GEN_534 = 4'h5 == csrs_8_Index ? tlb_5_ASID : _GEN_533;
  wire [9:0] _GEN_535 = 4'h6 == csrs_8_Index ? tlb_6_ASID : _GEN_534;
  wire [9:0] _GEN_536 = 4'h7 == csrs_8_Index ? tlb_7_ASID : _GEN_535;
  wire [9:0] _GEN_537 = 4'h8 == csrs_8_Index ? tlb_8_ASID : _GEN_536;
  wire [9:0] _GEN_538 = 4'h9 == csrs_8_Index ? tlb_9_ASID : _GEN_537;
  wire [9:0] _GEN_539 = 4'ha == csrs_8_Index ? tlb_10_ASID : _GEN_538;
  wire [9:0] _GEN_540 = 4'hb == csrs_8_Index ? tlb_11_ASID : _GEN_539;
  wire [9:0] _GEN_541 = 4'hc == csrs_8_Index ? tlb_12_ASID : _GEN_540;
  wire [9:0] _GEN_542 = 4'hd == csrs_8_Index ? tlb_13_ASID : _GEN_541;
  wire [9:0] _GEN_543 = 4'he == csrs_8_Index ? tlb_14_ASID : _GEN_542;
  wire [9:0] _GEN_544 = 4'hf == csrs_8_Index ? tlb_15_ASID : _GEN_543;
  wire [5:0] _GEN_545 = _GEN_320 ? _GEN_336 : 6'h0;
  wire [18:0] _GEN_546 = _GEN_320 ? _GEN_352 : 19'h0;
  wire [19:0] _GEN_547 = _GEN_320 ? _GEN_368 : 20'h0;
  wire  _GEN_548 = _GEN_320 & _GEN_384;
  wire [1:0] _GEN_549 = _GEN_320 ? _GEN_400 : 2'h0;
  wire [1:0] _GEN_550 = _GEN_320 ? _GEN_416 : 2'h0;
  wire  _GEN_551 = _GEN_320 & _GEN_432;
  wire  _GEN_552 = _GEN_320 & _GEN_448;
  wire [19:0] _GEN_553 = _GEN_320 ? _GEN_464 : 20'h0;
  wire [1:0] _GEN_555 = _GEN_320 ? _GEN_480 : 2'h0;
  wire [1:0] _GEN_556 = _GEN_320 ? _GEN_496 : 2'h0;
  wire  _GEN_557 = _GEN_320 & _GEN_512;
  wire  _GEN_558 = _GEN_320 & _GEN_528;
  wire [9:0] _GEN_559 = _GEN_320 ? _GEN_544 : 10'h0;
  wire [18:0] _GEN_560 = 4'h0 == csrs_8_Index ? csrs_9_VPPN : tlb_0_VPPN;
  wire [18:0] _GEN_561 = 4'h1 == csrs_8_Index ? csrs_9_VPPN : tlb_1_VPPN;
  wire [18:0] _GEN_562 = 4'h2 == csrs_8_Index ? csrs_9_VPPN : tlb_2_VPPN;
  wire [18:0] _GEN_563 = 4'h3 == csrs_8_Index ? csrs_9_VPPN : tlb_3_VPPN;
  wire [18:0] _GEN_564 = 4'h4 == csrs_8_Index ? csrs_9_VPPN : tlb_4_VPPN;
  wire [18:0] _GEN_565 = 4'h5 == csrs_8_Index ? csrs_9_VPPN : tlb_5_VPPN;
  wire [18:0] _GEN_566 = 4'h6 == csrs_8_Index ? csrs_9_VPPN : tlb_6_VPPN;
  wire [18:0] _GEN_567 = 4'h7 == csrs_8_Index ? csrs_9_VPPN : tlb_7_VPPN;
  wire [18:0] _GEN_568 = 4'h8 == csrs_8_Index ? csrs_9_VPPN : tlb_8_VPPN;
  wire [18:0] _GEN_569 = 4'h9 == csrs_8_Index ? csrs_9_VPPN : tlb_9_VPPN;
  wire [18:0] _GEN_570 = 4'ha == csrs_8_Index ? csrs_9_VPPN : tlb_10_VPPN;
  wire [18:0] _GEN_571 = 4'hb == csrs_8_Index ? csrs_9_VPPN : tlb_11_VPPN;
  wire [18:0] _GEN_572 = 4'hc == csrs_8_Index ? csrs_9_VPPN : tlb_12_VPPN;
  wire [18:0] _GEN_573 = 4'hd == csrs_8_Index ? csrs_9_VPPN : tlb_13_VPPN;
  wire [18:0] _GEN_574 = 4'he == csrs_8_Index ? csrs_9_VPPN : tlb_14_VPPN;
  wire [18:0] _GEN_575 = 4'hf == csrs_8_Index ? csrs_9_VPPN : tlb_15_VPPN;
  wire [5:0] _GEN_576 = 4'h0 == csrs_8_Index ? csrs_8_PS : tlb_0_PS;
  wire [5:0] _GEN_577 = 4'h1 == csrs_8_Index ? csrs_8_PS : tlb_1_PS;
  wire [5:0] _GEN_578 = 4'h2 == csrs_8_Index ? csrs_8_PS : tlb_2_PS;
  wire [5:0] _GEN_579 = 4'h3 == csrs_8_Index ? csrs_8_PS : tlb_3_PS;
  wire [5:0] _GEN_580 = 4'h4 == csrs_8_Index ? csrs_8_PS : tlb_4_PS;
  wire [5:0] _GEN_581 = 4'h5 == csrs_8_Index ? csrs_8_PS : tlb_5_PS;
  wire [5:0] _GEN_582 = 4'h6 == csrs_8_Index ? csrs_8_PS : tlb_6_PS;
  wire [5:0] _GEN_583 = 4'h7 == csrs_8_Index ? csrs_8_PS : tlb_7_PS;
  wire [5:0] _GEN_584 = 4'h8 == csrs_8_Index ? csrs_8_PS : tlb_8_PS;
  wire [5:0] _GEN_585 = 4'h9 == csrs_8_Index ? csrs_8_PS : tlb_9_PS;
  wire [5:0] _GEN_586 = 4'ha == csrs_8_Index ? csrs_8_PS : tlb_10_PS;
  wire [5:0] _GEN_587 = 4'hb == csrs_8_Index ? csrs_8_PS : tlb_11_PS;
  wire [5:0] _GEN_588 = 4'hc == csrs_8_Index ? csrs_8_PS : tlb_12_PS;
  wire [5:0] _GEN_589 = 4'hd == csrs_8_Index ? csrs_8_PS : tlb_13_PS;
  wire [5:0] _GEN_590 = 4'he == csrs_8_Index ? csrs_8_PS : tlb_14_PS;
  wire [5:0] _GEN_591 = 4'hf == csrs_8_Index ? csrs_8_PS : tlb_15_PS;
  wire  _GEN_592 = 4'h0 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_0_G;
  wire  _GEN_593 = 4'h1 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_1_G;
  wire  _GEN_594 = 4'h2 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_2_G;
  wire  _GEN_595 = 4'h3 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_3_G;
  wire  _GEN_596 = 4'h4 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_4_G;
  wire  _GEN_597 = 4'h5 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_5_G;
  wire  _GEN_598 = 4'h6 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_6_G;
  wire  _GEN_599 = 4'h7 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_7_G;
  wire  _GEN_600 = 4'h8 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_8_G;
  wire  _GEN_601 = 4'h9 == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_9_G;
  wire  _GEN_602 = 4'ha == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_10_G;
  wire  _GEN_603 = 4'hb == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_11_G;
  wire  _GEN_604 = 4'hc == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_12_G;
  wire  _GEN_605 = 4'hd == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_13_G;
  wire  _GEN_606 = 4'he == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_14_G;
  wire  _GEN_607 = 4'hf == csrs_8_Index ? csrs_10_G & csrs_11_G : tlb_15_G;
  wire [9:0] _GEN_608 = 4'h0 == csrs_8_Index ? asid_ASID : tlb_0_ASID;
  wire [9:0] _GEN_609 = 4'h1 == csrs_8_Index ? asid_ASID : tlb_1_ASID;
  wire [9:0] _GEN_610 = 4'h2 == csrs_8_Index ? asid_ASID : tlb_2_ASID;
  wire [9:0] _GEN_611 = 4'h3 == csrs_8_Index ? asid_ASID : tlb_3_ASID;
  wire [9:0] _GEN_612 = 4'h4 == csrs_8_Index ? asid_ASID : tlb_4_ASID;
  wire [9:0] _GEN_613 = 4'h5 == csrs_8_Index ? asid_ASID : tlb_5_ASID;
  wire [9:0] _GEN_614 = 4'h6 == csrs_8_Index ? asid_ASID : tlb_6_ASID;
  wire [9:0] _GEN_615 = 4'h7 == csrs_8_Index ? asid_ASID : tlb_7_ASID;
  wire [9:0] _GEN_616 = 4'h8 == csrs_8_Index ? asid_ASID : tlb_8_ASID;
  wire [9:0] _GEN_617 = 4'h9 == csrs_8_Index ? asid_ASID : tlb_9_ASID;
  wire [9:0] _GEN_618 = 4'ha == csrs_8_Index ? asid_ASID : tlb_10_ASID;
  wire [9:0] _GEN_619 = 4'hb == csrs_8_Index ? asid_ASID : tlb_11_ASID;
  wire [9:0] _GEN_620 = 4'hc == csrs_8_Index ? asid_ASID : tlb_12_ASID;
  wire [9:0] _GEN_621 = 4'hd == csrs_8_Index ? asid_ASID : tlb_13_ASID;
  wire [9:0] _GEN_622 = 4'he == csrs_8_Index ? asid_ASID : tlb_14_ASID;
  wire [9:0] _GEN_623 = 4'hf == csrs_8_Index ? asid_ASID : tlb_15_ASID;
  wire  _tlb_E_T = csrs_4_Ecode == 6'h3f;
  wire  _GEN_624 = 4'h0 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_0_E;
  wire  _GEN_625 = 4'h1 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_1_E;
  wire  _GEN_626 = 4'h2 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_2_E;
  wire  _GEN_627 = 4'h3 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_3_E;
  wire  _GEN_628 = 4'h4 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_4_E;
  wire  _GEN_629 = 4'h5 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_5_E;
  wire  _GEN_630 = 4'h6 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_6_E;
  wire  _GEN_631 = 4'h7 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_7_E;
  wire  _GEN_632 = 4'h8 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_8_E;
  wire  _GEN_633 = 4'h9 == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_9_E;
  wire  _GEN_634 = 4'ha == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_10_E;
  wire  _GEN_635 = 4'hb == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_11_E;
  wire  _GEN_636 = 4'hc == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_12_E;
  wire  _GEN_637 = 4'hd == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_13_E;
  wire  _GEN_638 = 4'he == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_14_E;
  wire  _GEN_639 = 4'hf == csrs_8_Index ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_15_E;
  wire [19:0] _GEN_640 = 4'h0 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_0_P0_PPN;
  wire [19:0] _GEN_641 = 4'h1 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_1_P0_PPN;
  wire [19:0] _GEN_642 = 4'h2 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_2_P0_PPN;
  wire [19:0] _GEN_643 = 4'h3 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_3_P0_PPN;
  wire [19:0] _GEN_644 = 4'h4 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_4_P0_PPN;
  wire [19:0] _GEN_645 = 4'h5 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_5_P0_PPN;
  wire [19:0] _GEN_646 = 4'h6 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_6_P0_PPN;
  wire [19:0] _GEN_647 = 4'h7 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_7_P0_PPN;
  wire [19:0] _GEN_648 = 4'h8 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_8_P0_PPN;
  wire [19:0] _GEN_649 = 4'h9 == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_9_P0_PPN;
  wire [19:0] _GEN_650 = 4'ha == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_10_P0_PPN;
  wire [19:0] _GEN_651 = 4'hb == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_11_P0_PPN;
  wire [19:0] _GEN_652 = 4'hc == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_12_P0_PPN;
  wire [19:0] _GEN_653 = 4'hd == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_13_P0_PPN;
  wire [19:0] _GEN_654 = 4'he == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_14_P0_PPN;
  wire [19:0] _GEN_655 = 4'hf == csrs_8_Index ? csrs_10_PPN[19:0] : tlb_15_P0_PPN;
  wire [1:0] _GEN_656 = 4'h0 == csrs_8_Index ? csrs_10_PLV : tlb_0_P0_PLV;
  wire [1:0] _GEN_657 = 4'h1 == csrs_8_Index ? csrs_10_PLV : tlb_1_P0_PLV;
  wire [1:0] _GEN_658 = 4'h2 == csrs_8_Index ? csrs_10_PLV : tlb_2_P0_PLV;
  wire [1:0] _GEN_659 = 4'h3 == csrs_8_Index ? csrs_10_PLV : tlb_3_P0_PLV;
  wire [1:0] _GEN_660 = 4'h4 == csrs_8_Index ? csrs_10_PLV : tlb_4_P0_PLV;
  wire [1:0] _GEN_661 = 4'h5 == csrs_8_Index ? csrs_10_PLV : tlb_5_P0_PLV;
  wire [1:0] _GEN_662 = 4'h6 == csrs_8_Index ? csrs_10_PLV : tlb_6_P0_PLV;
  wire [1:0] _GEN_663 = 4'h7 == csrs_8_Index ? csrs_10_PLV : tlb_7_P0_PLV;
  wire [1:0] _GEN_664 = 4'h8 == csrs_8_Index ? csrs_10_PLV : tlb_8_P0_PLV;
  wire [1:0] _GEN_665 = 4'h9 == csrs_8_Index ? csrs_10_PLV : tlb_9_P0_PLV;
  wire [1:0] _GEN_666 = 4'ha == csrs_8_Index ? csrs_10_PLV : tlb_10_P0_PLV;
  wire [1:0] _GEN_667 = 4'hb == csrs_8_Index ? csrs_10_PLV : tlb_11_P0_PLV;
  wire [1:0] _GEN_668 = 4'hc == csrs_8_Index ? csrs_10_PLV : tlb_12_P0_PLV;
  wire [1:0] _GEN_669 = 4'hd == csrs_8_Index ? csrs_10_PLV : tlb_13_P0_PLV;
  wire [1:0] _GEN_670 = 4'he == csrs_8_Index ? csrs_10_PLV : tlb_14_P0_PLV;
  wire [1:0] _GEN_671 = 4'hf == csrs_8_Index ? csrs_10_PLV : tlb_15_P0_PLV;
  wire [1:0] _GEN_672 = 4'h0 == csrs_8_Index ? csrs_10_MAT : tlb_0_P0_MAT;
  wire [1:0] _GEN_673 = 4'h1 == csrs_8_Index ? csrs_10_MAT : tlb_1_P0_MAT;
  wire [1:0] _GEN_674 = 4'h2 == csrs_8_Index ? csrs_10_MAT : tlb_2_P0_MAT;
  wire [1:0] _GEN_675 = 4'h3 == csrs_8_Index ? csrs_10_MAT : tlb_3_P0_MAT;
  wire [1:0] _GEN_676 = 4'h4 == csrs_8_Index ? csrs_10_MAT : tlb_4_P0_MAT;
  wire [1:0] _GEN_677 = 4'h5 == csrs_8_Index ? csrs_10_MAT : tlb_5_P0_MAT;
  wire [1:0] _GEN_678 = 4'h6 == csrs_8_Index ? csrs_10_MAT : tlb_6_P0_MAT;
  wire [1:0] _GEN_679 = 4'h7 == csrs_8_Index ? csrs_10_MAT : tlb_7_P0_MAT;
  wire [1:0] _GEN_680 = 4'h8 == csrs_8_Index ? csrs_10_MAT : tlb_8_P0_MAT;
  wire [1:0] _GEN_681 = 4'h9 == csrs_8_Index ? csrs_10_MAT : tlb_9_P0_MAT;
  wire [1:0] _GEN_682 = 4'ha == csrs_8_Index ? csrs_10_MAT : tlb_10_P0_MAT;
  wire [1:0] _GEN_683 = 4'hb == csrs_8_Index ? csrs_10_MAT : tlb_11_P0_MAT;
  wire [1:0] _GEN_684 = 4'hc == csrs_8_Index ? csrs_10_MAT : tlb_12_P0_MAT;
  wire [1:0] _GEN_685 = 4'hd == csrs_8_Index ? csrs_10_MAT : tlb_13_P0_MAT;
  wire [1:0] _GEN_686 = 4'he == csrs_8_Index ? csrs_10_MAT : tlb_14_P0_MAT;
  wire [1:0] _GEN_687 = 4'hf == csrs_8_Index ? csrs_10_MAT : tlb_15_P0_MAT;
  wire  _GEN_688 = 4'h0 == csrs_8_Index ? csrs_10_D : tlb_0_P0_D;
  wire  _GEN_689 = 4'h1 == csrs_8_Index ? csrs_10_D : tlb_1_P0_D;
  wire  _GEN_690 = 4'h2 == csrs_8_Index ? csrs_10_D : tlb_2_P0_D;
  wire  _GEN_691 = 4'h3 == csrs_8_Index ? csrs_10_D : tlb_3_P0_D;
  wire  _GEN_692 = 4'h4 == csrs_8_Index ? csrs_10_D : tlb_4_P0_D;
  wire  _GEN_693 = 4'h5 == csrs_8_Index ? csrs_10_D : tlb_5_P0_D;
  wire  _GEN_694 = 4'h6 == csrs_8_Index ? csrs_10_D : tlb_6_P0_D;
  wire  _GEN_695 = 4'h7 == csrs_8_Index ? csrs_10_D : tlb_7_P0_D;
  wire  _GEN_696 = 4'h8 == csrs_8_Index ? csrs_10_D : tlb_8_P0_D;
  wire  _GEN_697 = 4'h9 == csrs_8_Index ? csrs_10_D : tlb_9_P0_D;
  wire  _GEN_698 = 4'ha == csrs_8_Index ? csrs_10_D : tlb_10_P0_D;
  wire  _GEN_699 = 4'hb == csrs_8_Index ? csrs_10_D : tlb_11_P0_D;
  wire  _GEN_700 = 4'hc == csrs_8_Index ? csrs_10_D : tlb_12_P0_D;
  wire  _GEN_701 = 4'hd == csrs_8_Index ? csrs_10_D : tlb_13_P0_D;
  wire  _GEN_702 = 4'he == csrs_8_Index ? csrs_10_D : tlb_14_P0_D;
  wire  _GEN_703 = 4'hf == csrs_8_Index ? csrs_10_D : tlb_15_P0_D;
  wire  _GEN_704 = 4'h0 == csrs_8_Index ? csrs_10_V : tlb_0_P0_V;
  wire  _GEN_705 = 4'h1 == csrs_8_Index ? csrs_10_V : tlb_1_P0_V;
  wire  _GEN_706 = 4'h2 == csrs_8_Index ? csrs_10_V : tlb_2_P0_V;
  wire  _GEN_707 = 4'h3 == csrs_8_Index ? csrs_10_V : tlb_3_P0_V;
  wire  _GEN_708 = 4'h4 == csrs_8_Index ? csrs_10_V : tlb_4_P0_V;
  wire  _GEN_709 = 4'h5 == csrs_8_Index ? csrs_10_V : tlb_5_P0_V;
  wire  _GEN_710 = 4'h6 == csrs_8_Index ? csrs_10_V : tlb_6_P0_V;
  wire  _GEN_711 = 4'h7 == csrs_8_Index ? csrs_10_V : tlb_7_P0_V;
  wire  _GEN_712 = 4'h8 == csrs_8_Index ? csrs_10_V : tlb_8_P0_V;
  wire  _GEN_713 = 4'h9 == csrs_8_Index ? csrs_10_V : tlb_9_P0_V;
  wire  _GEN_714 = 4'ha == csrs_8_Index ? csrs_10_V : tlb_10_P0_V;
  wire  _GEN_715 = 4'hb == csrs_8_Index ? csrs_10_V : tlb_11_P0_V;
  wire  _GEN_716 = 4'hc == csrs_8_Index ? csrs_10_V : tlb_12_P0_V;
  wire  _GEN_717 = 4'hd == csrs_8_Index ? csrs_10_V : tlb_13_P0_V;
  wire  _GEN_718 = 4'he == csrs_8_Index ? csrs_10_V : tlb_14_P0_V;
  wire  _GEN_719 = 4'hf == csrs_8_Index ? csrs_10_V : tlb_15_P0_V;
  wire [19:0] _GEN_720 = 4'h0 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_0_P1_PPN;
  wire [19:0] _GEN_721 = 4'h1 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_1_P1_PPN;
  wire [19:0] _GEN_722 = 4'h2 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_2_P1_PPN;
  wire [19:0] _GEN_723 = 4'h3 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_3_P1_PPN;
  wire [19:0] _GEN_724 = 4'h4 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_4_P1_PPN;
  wire [19:0] _GEN_725 = 4'h5 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_5_P1_PPN;
  wire [19:0] _GEN_726 = 4'h6 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_6_P1_PPN;
  wire [19:0] _GEN_727 = 4'h7 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_7_P1_PPN;
  wire [19:0] _GEN_728 = 4'h8 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_8_P1_PPN;
  wire [19:0] _GEN_729 = 4'h9 == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_9_P1_PPN;
  wire [19:0] _GEN_730 = 4'ha == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_10_P1_PPN;
  wire [19:0] _GEN_731 = 4'hb == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_11_P1_PPN;
  wire [19:0] _GEN_732 = 4'hc == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_12_P1_PPN;
  wire [19:0] _GEN_733 = 4'hd == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_13_P1_PPN;
  wire [19:0] _GEN_734 = 4'he == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_14_P1_PPN;
  wire [19:0] _GEN_735 = 4'hf == csrs_8_Index ? csrs_11_PPN[19:0] : tlb_15_P1_PPN;
  wire [1:0] _GEN_736 = 4'h0 == csrs_8_Index ? csrs_11_PLV : tlb_0_P1_PLV;
  wire [1:0] _GEN_737 = 4'h1 == csrs_8_Index ? csrs_11_PLV : tlb_1_P1_PLV;
  wire [1:0] _GEN_738 = 4'h2 == csrs_8_Index ? csrs_11_PLV : tlb_2_P1_PLV;
  wire [1:0] _GEN_739 = 4'h3 == csrs_8_Index ? csrs_11_PLV : tlb_3_P1_PLV;
  wire [1:0] _GEN_740 = 4'h4 == csrs_8_Index ? csrs_11_PLV : tlb_4_P1_PLV;
  wire [1:0] _GEN_741 = 4'h5 == csrs_8_Index ? csrs_11_PLV : tlb_5_P1_PLV;
  wire [1:0] _GEN_742 = 4'h6 == csrs_8_Index ? csrs_11_PLV : tlb_6_P1_PLV;
  wire [1:0] _GEN_743 = 4'h7 == csrs_8_Index ? csrs_11_PLV : tlb_7_P1_PLV;
  wire [1:0] _GEN_744 = 4'h8 == csrs_8_Index ? csrs_11_PLV : tlb_8_P1_PLV;
  wire [1:0] _GEN_745 = 4'h9 == csrs_8_Index ? csrs_11_PLV : tlb_9_P1_PLV;
  wire [1:0] _GEN_746 = 4'ha == csrs_8_Index ? csrs_11_PLV : tlb_10_P1_PLV;
  wire [1:0] _GEN_747 = 4'hb == csrs_8_Index ? csrs_11_PLV : tlb_11_P1_PLV;
  wire [1:0] _GEN_748 = 4'hc == csrs_8_Index ? csrs_11_PLV : tlb_12_P1_PLV;
  wire [1:0] _GEN_749 = 4'hd == csrs_8_Index ? csrs_11_PLV : tlb_13_P1_PLV;
  wire [1:0] _GEN_750 = 4'he == csrs_8_Index ? csrs_11_PLV : tlb_14_P1_PLV;
  wire [1:0] _GEN_751 = 4'hf == csrs_8_Index ? csrs_11_PLV : tlb_15_P1_PLV;
  wire [1:0] _GEN_752 = 4'h0 == csrs_8_Index ? csrs_11_MAT : tlb_0_P1_MAT;
  wire [1:0] _GEN_753 = 4'h1 == csrs_8_Index ? csrs_11_MAT : tlb_1_P1_MAT;
  wire [1:0] _GEN_754 = 4'h2 == csrs_8_Index ? csrs_11_MAT : tlb_2_P1_MAT;
  wire [1:0] _GEN_755 = 4'h3 == csrs_8_Index ? csrs_11_MAT : tlb_3_P1_MAT;
  wire [1:0] _GEN_756 = 4'h4 == csrs_8_Index ? csrs_11_MAT : tlb_4_P1_MAT;
  wire [1:0] _GEN_757 = 4'h5 == csrs_8_Index ? csrs_11_MAT : tlb_5_P1_MAT;
  wire [1:0] _GEN_758 = 4'h6 == csrs_8_Index ? csrs_11_MAT : tlb_6_P1_MAT;
  wire [1:0] _GEN_759 = 4'h7 == csrs_8_Index ? csrs_11_MAT : tlb_7_P1_MAT;
  wire [1:0] _GEN_760 = 4'h8 == csrs_8_Index ? csrs_11_MAT : tlb_8_P1_MAT;
  wire [1:0] _GEN_761 = 4'h9 == csrs_8_Index ? csrs_11_MAT : tlb_9_P1_MAT;
  wire [1:0] _GEN_762 = 4'ha == csrs_8_Index ? csrs_11_MAT : tlb_10_P1_MAT;
  wire [1:0] _GEN_763 = 4'hb == csrs_8_Index ? csrs_11_MAT : tlb_11_P1_MAT;
  wire [1:0] _GEN_764 = 4'hc == csrs_8_Index ? csrs_11_MAT : tlb_12_P1_MAT;
  wire [1:0] _GEN_765 = 4'hd == csrs_8_Index ? csrs_11_MAT : tlb_13_P1_MAT;
  wire [1:0] _GEN_766 = 4'he == csrs_8_Index ? csrs_11_MAT : tlb_14_P1_MAT;
  wire [1:0] _GEN_767 = 4'hf == csrs_8_Index ? csrs_11_MAT : tlb_15_P1_MAT;
  wire  _GEN_768 = 4'h0 == csrs_8_Index ? csrs_11_D : tlb_0_P1_D;
  wire  _GEN_769 = 4'h1 == csrs_8_Index ? csrs_11_D : tlb_1_P1_D;
  wire  _GEN_770 = 4'h2 == csrs_8_Index ? csrs_11_D : tlb_2_P1_D;
  wire  _GEN_771 = 4'h3 == csrs_8_Index ? csrs_11_D : tlb_3_P1_D;
  wire  _GEN_772 = 4'h4 == csrs_8_Index ? csrs_11_D : tlb_4_P1_D;
  wire  _GEN_773 = 4'h5 == csrs_8_Index ? csrs_11_D : tlb_5_P1_D;
  wire  _GEN_774 = 4'h6 == csrs_8_Index ? csrs_11_D : tlb_6_P1_D;
  wire  _GEN_775 = 4'h7 == csrs_8_Index ? csrs_11_D : tlb_7_P1_D;
  wire  _GEN_776 = 4'h8 == csrs_8_Index ? csrs_11_D : tlb_8_P1_D;
  wire  _GEN_777 = 4'h9 == csrs_8_Index ? csrs_11_D : tlb_9_P1_D;
  wire  _GEN_778 = 4'ha == csrs_8_Index ? csrs_11_D : tlb_10_P1_D;
  wire  _GEN_779 = 4'hb == csrs_8_Index ? csrs_11_D : tlb_11_P1_D;
  wire  _GEN_780 = 4'hc == csrs_8_Index ? csrs_11_D : tlb_12_P1_D;
  wire  _GEN_781 = 4'hd == csrs_8_Index ? csrs_11_D : tlb_13_P1_D;
  wire  _GEN_782 = 4'he == csrs_8_Index ? csrs_11_D : tlb_14_P1_D;
  wire  _GEN_783 = 4'hf == csrs_8_Index ? csrs_11_D : tlb_15_P1_D;
  wire  _GEN_784 = 4'h0 == csrs_8_Index ? csrs_11_V : tlb_0_P1_V;
  wire  _GEN_785 = 4'h1 == csrs_8_Index ? csrs_11_V : tlb_1_P1_V;
  wire  _GEN_786 = 4'h2 == csrs_8_Index ? csrs_11_V : tlb_2_P1_V;
  wire  _GEN_787 = 4'h3 == csrs_8_Index ? csrs_11_V : tlb_3_P1_V;
  wire  _GEN_788 = 4'h4 == csrs_8_Index ? csrs_11_V : tlb_4_P1_V;
  wire  _GEN_789 = 4'h5 == csrs_8_Index ? csrs_11_V : tlb_5_P1_V;
  wire  _GEN_790 = 4'h6 == csrs_8_Index ? csrs_11_V : tlb_6_P1_V;
  wire  _GEN_791 = 4'h7 == csrs_8_Index ? csrs_11_V : tlb_7_P1_V;
  wire  _GEN_792 = 4'h8 == csrs_8_Index ? csrs_11_V : tlb_8_P1_V;
  wire  _GEN_793 = 4'h9 == csrs_8_Index ? csrs_11_V : tlb_9_P1_V;
  wire  _GEN_794 = 4'ha == csrs_8_Index ? csrs_11_V : tlb_10_P1_V;
  wire  _GEN_795 = 4'hb == csrs_8_Index ? csrs_11_V : tlb_11_P1_V;
  wire  _GEN_796 = 4'hc == csrs_8_Index ? csrs_11_V : tlb_12_P1_V;
  wire  _GEN_797 = 4'hd == csrs_8_Index ? csrs_11_V : tlb_13_P1_V;
  wire  _GEN_798 = 4'he == csrs_8_Index ? csrs_11_V : tlb_14_P1_V;
  wire  _GEN_799 = 4'hf == csrs_8_Index ? csrs_11_V : tlb_15_P1_V;
  wire [18:0] _GEN_800 = 4'h0 == timer[3:0] ? csrs_9_VPPN : tlb_0_VPPN;
  wire [18:0] _GEN_801 = 4'h1 == timer[3:0] ? csrs_9_VPPN : tlb_1_VPPN;
  wire [18:0] _GEN_802 = 4'h2 == timer[3:0] ? csrs_9_VPPN : tlb_2_VPPN;
  wire [18:0] _GEN_803 = 4'h3 == timer[3:0] ? csrs_9_VPPN : tlb_3_VPPN;
  wire [18:0] _GEN_804 = 4'h4 == timer[3:0] ? csrs_9_VPPN : tlb_4_VPPN;
  wire [18:0] _GEN_805 = 4'h5 == timer[3:0] ? csrs_9_VPPN : tlb_5_VPPN;
  wire [18:0] _GEN_806 = 4'h6 == timer[3:0] ? csrs_9_VPPN : tlb_6_VPPN;
  wire [18:0] _GEN_807 = 4'h7 == timer[3:0] ? csrs_9_VPPN : tlb_7_VPPN;
  wire [18:0] _GEN_808 = 4'h8 == timer[3:0] ? csrs_9_VPPN : tlb_8_VPPN;
  wire [18:0] _GEN_809 = 4'h9 == timer[3:0] ? csrs_9_VPPN : tlb_9_VPPN;
  wire [18:0] _GEN_810 = 4'ha == timer[3:0] ? csrs_9_VPPN : tlb_10_VPPN;
  wire [18:0] _GEN_811 = 4'hb == timer[3:0] ? csrs_9_VPPN : tlb_11_VPPN;
  wire [18:0] _GEN_812 = 4'hc == timer[3:0] ? csrs_9_VPPN : tlb_12_VPPN;
  wire [18:0] _GEN_813 = 4'hd == timer[3:0] ? csrs_9_VPPN : tlb_13_VPPN;
  wire [18:0] _GEN_814 = 4'he == timer[3:0] ? csrs_9_VPPN : tlb_14_VPPN;
  wire [18:0] _GEN_815 = 4'hf == timer[3:0] ? csrs_9_VPPN : tlb_15_VPPN;
  wire [5:0] _GEN_816 = 4'h0 == timer[3:0] ? csrs_8_PS : tlb_0_PS;
  wire [5:0] _GEN_817 = 4'h1 == timer[3:0] ? csrs_8_PS : tlb_1_PS;
  wire [5:0] _GEN_818 = 4'h2 == timer[3:0] ? csrs_8_PS : tlb_2_PS;
  wire [5:0] _GEN_819 = 4'h3 == timer[3:0] ? csrs_8_PS : tlb_3_PS;
  wire [5:0] _GEN_820 = 4'h4 == timer[3:0] ? csrs_8_PS : tlb_4_PS;
  wire [5:0] _GEN_821 = 4'h5 == timer[3:0] ? csrs_8_PS : tlb_5_PS;
  wire [5:0] _GEN_822 = 4'h6 == timer[3:0] ? csrs_8_PS : tlb_6_PS;
  wire [5:0] _GEN_823 = 4'h7 == timer[3:0] ? csrs_8_PS : tlb_7_PS;
  wire [5:0] _GEN_824 = 4'h8 == timer[3:0] ? csrs_8_PS : tlb_8_PS;
  wire [5:0] _GEN_825 = 4'h9 == timer[3:0] ? csrs_8_PS : tlb_9_PS;
  wire [5:0] _GEN_826 = 4'ha == timer[3:0] ? csrs_8_PS : tlb_10_PS;
  wire [5:0] _GEN_827 = 4'hb == timer[3:0] ? csrs_8_PS : tlb_11_PS;
  wire [5:0] _GEN_828 = 4'hc == timer[3:0] ? csrs_8_PS : tlb_12_PS;
  wire [5:0] _GEN_829 = 4'hd == timer[3:0] ? csrs_8_PS : tlb_13_PS;
  wire [5:0] _GEN_830 = 4'he == timer[3:0] ? csrs_8_PS : tlb_14_PS;
  wire [5:0] _GEN_831 = 4'hf == timer[3:0] ? csrs_8_PS : tlb_15_PS;
  wire  _GEN_832 = 4'h0 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_0_G;
  wire  _GEN_833 = 4'h1 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_1_G;
  wire  _GEN_834 = 4'h2 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_2_G;
  wire  _GEN_835 = 4'h3 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_3_G;
  wire  _GEN_836 = 4'h4 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_4_G;
  wire  _GEN_837 = 4'h5 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_5_G;
  wire  _GEN_838 = 4'h6 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_6_G;
  wire  _GEN_839 = 4'h7 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_7_G;
  wire  _GEN_840 = 4'h8 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_8_G;
  wire  _GEN_841 = 4'h9 == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_9_G;
  wire  _GEN_842 = 4'ha == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_10_G;
  wire  _GEN_843 = 4'hb == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_11_G;
  wire  _GEN_844 = 4'hc == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_12_G;
  wire  _GEN_845 = 4'hd == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_13_G;
  wire  _GEN_846 = 4'he == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_14_G;
  wire  _GEN_847 = 4'hf == timer[3:0] ? csrs_10_G & csrs_11_G : tlb_15_G;
  wire [9:0] _GEN_848 = 4'h0 == timer[3:0] ? asid_ASID : tlb_0_ASID;
  wire [9:0] _GEN_849 = 4'h1 == timer[3:0] ? asid_ASID : tlb_1_ASID;
  wire [9:0] _GEN_850 = 4'h2 == timer[3:0] ? asid_ASID : tlb_2_ASID;
  wire [9:0] _GEN_851 = 4'h3 == timer[3:0] ? asid_ASID : tlb_3_ASID;
  wire [9:0] _GEN_852 = 4'h4 == timer[3:0] ? asid_ASID : tlb_4_ASID;
  wire [9:0] _GEN_853 = 4'h5 == timer[3:0] ? asid_ASID : tlb_5_ASID;
  wire [9:0] _GEN_854 = 4'h6 == timer[3:0] ? asid_ASID : tlb_6_ASID;
  wire [9:0] _GEN_855 = 4'h7 == timer[3:0] ? asid_ASID : tlb_7_ASID;
  wire [9:0] _GEN_856 = 4'h8 == timer[3:0] ? asid_ASID : tlb_8_ASID;
  wire [9:0] _GEN_857 = 4'h9 == timer[3:0] ? asid_ASID : tlb_9_ASID;
  wire [9:0] _GEN_858 = 4'ha == timer[3:0] ? asid_ASID : tlb_10_ASID;
  wire [9:0] _GEN_859 = 4'hb == timer[3:0] ? asid_ASID : tlb_11_ASID;
  wire [9:0] _GEN_860 = 4'hc == timer[3:0] ? asid_ASID : tlb_12_ASID;
  wire [9:0] _GEN_861 = 4'hd == timer[3:0] ? asid_ASID : tlb_13_ASID;
  wire [9:0] _GEN_862 = 4'he == timer[3:0] ? asid_ASID : tlb_14_ASID;
  wire [9:0] _GEN_863 = 4'hf == timer[3:0] ? asid_ASID : tlb_15_ASID;
  wire  _GEN_864 = 4'h0 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_0_E;
  wire  _GEN_865 = 4'h1 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_1_E;
  wire  _GEN_866 = 4'h2 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_2_E;
  wire  _GEN_867 = 4'h3 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_3_E;
  wire  _GEN_868 = 4'h4 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_4_E;
  wire  _GEN_869 = 4'h5 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_5_E;
  wire  _GEN_870 = 4'h6 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_6_E;
  wire  _GEN_871 = 4'h7 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_7_E;
  wire  _GEN_872 = 4'h8 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_8_E;
  wire  _GEN_873 = 4'h9 == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_9_E;
  wire  _GEN_874 = 4'ha == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_10_E;
  wire  _GEN_875 = 4'hb == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_11_E;
  wire  _GEN_876 = 4'hc == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_12_E;
  wire  _GEN_877 = 4'hd == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_13_E;
  wire  _GEN_878 = 4'he == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_14_E;
  wire  _GEN_879 = 4'hf == timer[3:0] ? csrs_4_Ecode == 6'h3f | ~csrs_8_NE : tlb_15_E;
  wire [19:0] _GEN_880 = 4'h0 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_0_P0_PPN;
  wire [19:0] _GEN_881 = 4'h1 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_1_P0_PPN;
  wire [19:0] _GEN_882 = 4'h2 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_2_P0_PPN;
  wire [19:0] _GEN_883 = 4'h3 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_3_P0_PPN;
  wire [19:0] _GEN_884 = 4'h4 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_4_P0_PPN;
  wire [19:0] _GEN_885 = 4'h5 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_5_P0_PPN;
  wire [19:0] _GEN_886 = 4'h6 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_6_P0_PPN;
  wire [19:0] _GEN_887 = 4'h7 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_7_P0_PPN;
  wire [19:0] _GEN_888 = 4'h8 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_8_P0_PPN;
  wire [19:0] _GEN_889 = 4'h9 == timer[3:0] ? csrs_10_PPN[19:0] : tlb_9_P0_PPN;
  wire [19:0] _GEN_890 = 4'ha == timer[3:0] ? csrs_10_PPN[19:0] : tlb_10_P0_PPN;
  wire [19:0] _GEN_891 = 4'hb == timer[3:0] ? csrs_10_PPN[19:0] : tlb_11_P0_PPN;
  wire [19:0] _GEN_892 = 4'hc == timer[3:0] ? csrs_10_PPN[19:0] : tlb_12_P0_PPN;
  wire [19:0] _GEN_893 = 4'hd == timer[3:0] ? csrs_10_PPN[19:0] : tlb_13_P0_PPN;
  wire [19:0] _GEN_894 = 4'he == timer[3:0] ? csrs_10_PPN[19:0] : tlb_14_P0_PPN;
  wire [19:0] _GEN_895 = 4'hf == timer[3:0] ? csrs_10_PPN[19:0] : tlb_15_P0_PPN;
  wire [1:0] _GEN_896 = 4'h0 == timer[3:0] ? csrs_10_PLV : tlb_0_P0_PLV;
  wire [1:0] _GEN_897 = 4'h1 == timer[3:0] ? csrs_10_PLV : tlb_1_P0_PLV;
  wire [1:0] _GEN_898 = 4'h2 == timer[3:0] ? csrs_10_PLV : tlb_2_P0_PLV;
  wire [1:0] _GEN_899 = 4'h3 == timer[3:0] ? csrs_10_PLV : tlb_3_P0_PLV;
  wire [1:0] _GEN_900 = 4'h4 == timer[3:0] ? csrs_10_PLV : tlb_4_P0_PLV;
  wire [1:0] _GEN_901 = 4'h5 == timer[3:0] ? csrs_10_PLV : tlb_5_P0_PLV;
  wire [1:0] _GEN_902 = 4'h6 == timer[3:0] ? csrs_10_PLV : tlb_6_P0_PLV;
  wire [1:0] _GEN_903 = 4'h7 == timer[3:0] ? csrs_10_PLV : tlb_7_P0_PLV;
  wire [1:0] _GEN_904 = 4'h8 == timer[3:0] ? csrs_10_PLV : tlb_8_P0_PLV;
  wire [1:0] _GEN_905 = 4'h9 == timer[3:0] ? csrs_10_PLV : tlb_9_P0_PLV;
  wire [1:0] _GEN_906 = 4'ha == timer[3:0] ? csrs_10_PLV : tlb_10_P0_PLV;
  wire [1:0] _GEN_907 = 4'hb == timer[3:0] ? csrs_10_PLV : tlb_11_P0_PLV;
  wire [1:0] _GEN_908 = 4'hc == timer[3:0] ? csrs_10_PLV : tlb_12_P0_PLV;
  wire [1:0] _GEN_909 = 4'hd == timer[3:0] ? csrs_10_PLV : tlb_13_P0_PLV;
  wire [1:0] _GEN_910 = 4'he == timer[3:0] ? csrs_10_PLV : tlb_14_P0_PLV;
  wire [1:0] _GEN_911 = 4'hf == timer[3:0] ? csrs_10_PLV : tlb_15_P0_PLV;
  wire [1:0] _GEN_912 = 4'h0 == timer[3:0] ? csrs_10_MAT : tlb_0_P0_MAT;
  wire [1:0] _GEN_913 = 4'h1 == timer[3:0] ? csrs_10_MAT : tlb_1_P0_MAT;
  wire [1:0] _GEN_914 = 4'h2 == timer[3:0] ? csrs_10_MAT : tlb_2_P0_MAT;
  wire [1:0] _GEN_915 = 4'h3 == timer[3:0] ? csrs_10_MAT : tlb_3_P0_MAT;
  wire [1:0] _GEN_916 = 4'h4 == timer[3:0] ? csrs_10_MAT : tlb_4_P0_MAT;
  wire [1:0] _GEN_917 = 4'h5 == timer[3:0] ? csrs_10_MAT : tlb_5_P0_MAT;
  wire [1:0] _GEN_918 = 4'h6 == timer[3:0] ? csrs_10_MAT : tlb_6_P0_MAT;
  wire [1:0] _GEN_919 = 4'h7 == timer[3:0] ? csrs_10_MAT : tlb_7_P0_MAT;
  wire [1:0] _GEN_920 = 4'h8 == timer[3:0] ? csrs_10_MAT : tlb_8_P0_MAT;
  wire [1:0] _GEN_921 = 4'h9 == timer[3:0] ? csrs_10_MAT : tlb_9_P0_MAT;
  wire [1:0] _GEN_922 = 4'ha == timer[3:0] ? csrs_10_MAT : tlb_10_P0_MAT;
  wire [1:0] _GEN_923 = 4'hb == timer[3:0] ? csrs_10_MAT : tlb_11_P0_MAT;
  wire [1:0] _GEN_924 = 4'hc == timer[3:0] ? csrs_10_MAT : tlb_12_P0_MAT;
  wire [1:0] _GEN_925 = 4'hd == timer[3:0] ? csrs_10_MAT : tlb_13_P0_MAT;
  wire [1:0] _GEN_926 = 4'he == timer[3:0] ? csrs_10_MAT : tlb_14_P0_MAT;
  wire [1:0] _GEN_927 = 4'hf == timer[3:0] ? csrs_10_MAT : tlb_15_P0_MAT;
  wire  _GEN_928 = 4'h0 == timer[3:0] ? csrs_10_D : tlb_0_P0_D;
  wire  _GEN_929 = 4'h1 == timer[3:0] ? csrs_10_D : tlb_1_P0_D;
  wire  _GEN_930 = 4'h2 == timer[3:0] ? csrs_10_D : tlb_2_P0_D;
  wire  _GEN_931 = 4'h3 == timer[3:0] ? csrs_10_D : tlb_3_P0_D;
  wire  _GEN_932 = 4'h4 == timer[3:0] ? csrs_10_D : tlb_4_P0_D;
  wire  _GEN_933 = 4'h5 == timer[3:0] ? csrs_10_D : tlb_5_P0_D;
  wire  _GEN_934 = 4'h6 == timer[3:0] ? csrs_10_D : tlb_6_P0_D;
  wire  _GEN_935 = 4'h7 == timer[3:0] ? csrs_10_D : tlb_7_P0_D;
  wire  _GEN_936 = 4'h8 == timer[3:0] ? csrs_10_D : tlb_8_P0_D;
  wire  _GEN_937 = 4'h9 == timer[3:0] ? csrs_10_D : tlb_9_P0_D;
  wire  _GEN_938 = 4'ha == timer[3:0] ? csrs_10_D : tlb_10_P0_D;
  wire  _GEN_939 = 4'hb == timer[3:0] ? csrs_10_D : tlb_11_P0_D;
  wire  _GEN_940 = 4'hc == timer[3:0] ? csrs_10_D : tlb_12_P0_D;
  wire  _GEN_941 = 4'hd == timer[3:0] ? csrs_10_D : tlb_13_P0_D;
  wire  _GEN_942 = 4'he == timer[3:0] ? csrs_10_D : tlb_14_P0_D;
  wire  _GEN_943 = 4'hf == timer[3:0] ? csrs_10_D : tlb_15_P0_D;
  wire  _GEN_944 = 4'h0 == timer[3:0] ? csrs_10_V : tlb_0_P0_V;
  wire  _GEN_945 = 4'h1 == timer[3:0] ? csrs_10_V : tlb_1_P0_V;
  wire  _GEN_946 = 4'h2 == timer[3:0] ? csrs_10_V : tlb_2_P0_V;
  wire  _GEN_947 = 4'h3 == timer[3:0] ? csrs_10_V : tlb_3_P0_V;
  wire  _GEN_948 = 4'h4 == timer[3:0] ? csrs_10_V : tlb_4_P0_V;
  wire  _GEN_949 = 4'h5 == timer[3:0] ? csrs_10_V : tlb_5_P0_V;
  wire  _GEN_950 = 4'h6 == timer[3:0] ? csrs_10_V : tlb_6_P0_V;
  wire  _GEN_951 = 4'h7 == timer[3:0] ? csrs_10_V : tlb_7_P0_V;
  wire  _GEN_952 = 4'h8 == timer[3:0] ? csrs_10_V : tlb_8_P0_V;
  wire  _GEN_953 = 4'h9 == timer[3:0] ? csrs_10_V : tlb_9_P0_V;
  wire  _GEN_954 = 4'ha == timer[3:0] ? csrs_10_V : tlb_10_P0_V;
  wire  _GEN_955 = 4'hb == timer[3:0] ? csrs_10_V : tlb_11_P0_V;
  wire  _GEN_956 = 4'hc == timer[3:0] ? csrs_10_V : tlb_12_P0_V;
  wire  _GEN_957 = 4'hd == timer[3:0] ? csrs_10_V : tlb_13_P0_V;
  wire  _GEN_958 = 4'he == timer[3:0] ? csrs_10_V : tlb_14_P0_V;
  wire  _GEN_959 = 4'hf == timer[3:0] ? csrs_10_V : tlb_15_P0_V;
  wire [19:0] _GEN_960 = 4'h0 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_0_P1_PPN;
  wire [19:0] _GEN_961 = 4'h1 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_1_P1_PPN;
  wire [19:0] _GEN_962 = 4'h2 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_2_P1_PPN;
  wire [19:0] _GEN_963 = 4'h3 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_3_P1_PPN;
  wire [19:0] _GEN_964 = 4'h4 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_4_P1_PPN;
  wire [19:0] _GEN_965 = 4'h5 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_5_P1_PPN;
  wire [19:0] _GEN_966 = 4'h6 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_6_P1_PPN;
  wire [19:0] _GEN_967 = 4'h7 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_7_P1_PPN;
  wire [19:0] _GEN_968 = 4'h8 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_8_P1_PPN;
  wire [19:0] _GEN_969 = 4'h9 == timer[3:0] ? csrs_11_PPN[19:0] : tlb_9_P1_PPN;
  wire [19:0] _GEN_970 = 4'ha == timer[3:0] ? csrs_11_PPN[19:0] : tlb_10_P1_PPN;
  wire [19:0] _GEN_971 = 4'hb == timer[3:0] ? csrs_11_PPN[19:0] : tlb_11_P1_PPN;
  wire [19:0] _GEN_972 = 4'hc == timer[3:0] ? csrs_11_PPN[19:0] : tlb_12_P1_PPN;
  wire [19:0] _GEN_973 = 4'hd == timer[3:0] ? csrs_11_PPN[19:0] : tlb_13_P1_PPN;
  wire [19:0] _GEN_974 = 4'he == timer[3:0] ? csrs_11_PPN[19:0] : tlb_14_P1_PPN;
  wire [19:0] _GEN_975 = 4'hf == timer[3:0] ? csrs_11_PPN[19:0] : tlb_15_P1_PPN;
  wire [1:0] _GEN_976 = 4'h0 == timer[3:0] ? csrs_11_PLV : tlb_0_P1_PLV;
  wire [1:0] _GEN_977 = 4'h1 == timer[3:0] ? csrs_11_PLV : tlb_1_P1_PLV;
  wire [1:0] _GEN_978 = 4'h2 == timer[3:0] ? csrs_11_PLV : tlb_2_P1_PLV;
  wire [1:0] _GEN_979 = 4'h3 == timer[3:0] ? csrs_11_PLV : tlb_3_P1_PLV;
  wire [1:0] _GEN_980 = 4'h4 == timer[3:0] ? csrs_11_PLV : tlb_4_P1_PLV;
  wire [1:0] _GEN_981 = 4'h5 == timer[3:0] ? csrs_11_PLV : tlb_5_P1_PLV;
  wire [1:0] _GEN_982 = 4'h6 == timer[3:0] ? csrs_11_PLV : tlb_6_P1_PLV;
  wire [1:0] _GEN_983 = 4'h7 == timer[3:0] ? csrs_11_PLV : tlb_7_P1_PLV;
  wire [1:0] _GEN_984 = 4'h8 == timer[3:0] ? csrs_11_PLV : tlb_8_P1_PLV;
  wire [1:0] _GEN_985 = 4'h9 == timer[3:0] ? csrs_11_PLV : tlb_9_P1_PLV;
  wire [1:0] _GEN_986 = 4'ha == timer[3:0] ? csrs_11_PLV : tlb_10_P1_PLV;
  wire [1:0] _GEN_987 = 4'hb == timer[3:0] ? csrs_11_PLV : tlb_11_P1_PLV;
  wire [1:0] _GEN_988 = 4'hc == timer[3:0] ? csrs_11_PLV : tlb_12_P1_PLV;
  wire [1:0] _GEN_989 = 4'hd == timer[3:0] ? csrs_11_PLV : tlb_13_P1_PLV;
  wire [1:0] _GEN_990 = 4'he == timer[3:0] ? csrs_11_PLV : tlb_14_P1_PLV;
  wire [1:0] _GEN_991 = 4'hf == timer[3:0] ? csrs_11_PLV : tlb_15_P1_PLV;
  wire [1:0] _GEN_992 = 4'h0 == timer[3:0] ? csrs_11_MAT : tlb_0_P1_MAT;
  wire [1:0] _GEN_993 = 4'h1 == timer[3:0] ? csrs_11_MAT : tlb_1_P1_MAT;
  wire [1:0] _GEN_994 = 4'h2 == timer[3:0] ? csrs_11_MAT : tlb_2_P1_MAT;
  wire [1:0] _GEN_995 = 4'h3 == timer[3:0] ? csrs_11_MAT : tlb_3_P1_MAT;
  wire [1:0] _GEN_996 = 4'h4 == timer[3:0] ? csrs_11_MAT : tlb_4_P1_MAT;
  wire [1:0] _GEN_997 = 4'h5 == timer[3:0] ? csrs_11_MAT : tlb_5_P1_MAT;
  wire [1:0] _GEN_998 = 4'h6 == timer[3:0] ? csrs_11_MAT : tlb_6_P1_MAT;
  wire [1:0] _GEN_999 = 4'h7 == timer[3:0] ? csrs_11_MAT : tlb_7_P1_MAT;
  wire [1:0] _GEN_1000 = 4'h8 == timer[3:0] ? csrs_11_MAT : tlb_8_P1_MAT;
  wire [1:0] _GEN_1001 = 4'h9 == timer[3:0] ? csrs_11_MAT : tlb_9_P1_MAT;
  wire [1:0] _GEN_1002 = 4'ha == timer[3:0] ? csrs_11_MAT : tlb_10_P1_MAT;
  wire [1:0] _GEN_1003 = 4'hb == timer[3:0] ? csrs_11_MAT : tlb_11_P1_MAT;
  wire [1:0] _GEN_1004 = 4'hc == timer[3:0] ? csrs_11_MAT : tlb_12_P1_MAT;
  wire [1:0] _GEN_1005 = 4'hd == timer[3:0] ? csrs_11_MAT : tlb_13_P1_MAT;
  wire [1:0] _GEN_1006 = 4'he == timer[3:0] ? csrs_11_MAT : tlb_14_P1_MAT;
  wire [1:0] _GEN_1007 = 4'hf == timer[3:0] ? csrs_11_MAT : tlb_15_P1_MAT;
  wire  _GEN_1008 = 4'h0 == timer[3:0] ? csrs_11_D : tlb_0_P1_D;
  wire  _GEN_1009 = 4'h1 == timer[3:0] ? csrs_11_D : tlb_1_P1_D;
  wire  _GEN_1010 = 4'h2 == timer[3:0] ? csrs_11_D : tlb_2_P1_D;
  wire  _GEN_1011 = 4'h3 == timer[3:0] ? csrs_11_D : tlb_3_P1_D;
  wire  _GEN_1012 = 4'h4 == timer[3:0] ? csrs_11_D : tlb_4_P1_D;
  wire  _GEN_1013 = 4'h5 == timer[3:0] ? csrs_11_D : tlb_5_P1_D;
  wire  _GEN_1014 = 4'h6 == timer[3:0] ? csrs_11_D : tlb_6_P1_D;
  wire  _GEN_1015 = 4'h7 == timer[3:0] ? csrs_11_D : tlb_7_P1_D;
  wire  _GEN_1016 = 4'h8 == timer[3:0] ? csrs_11_D : tlb_8_P1_D;
  wire  _GEN_1017 = 4'h9 == timer[3:0] ? csrs_11_D : tlb_9_P1_D;
  wire  _GEN_1018 = 4'ha == timer[3:0] ? csrs_11_D : tlb_10_P1_D;
  wire  _GEN_1019 = 4'hb == timer[3:0] ? csrs_11_D : tlb_11_P1_D;
  wire  _GEN_1020 = 4'hc == timer[3:0] ? csrs_11_D : tlb_12_P1_D;
  wire  _GEN_1021 = 4'hd == timer[3:0] ? csrs_11_D : tlb_13_P1_D;
  wire  _GEN_1022 = 4'he == timer[3:0] ? csrs_11_D : tlb_14_P1_D;
  wire  _GEN_1023 = 4'hf == timer[3:0] ? csrs_11_D : tlb_15_P1_D;
  wire  _GEN_1024 = 4'h0 == timer[3:0] ? csrs_11_V : tlb_0_P1_V;
  wire  _GEN_1025 = 4'h1 == timer[3:0] ? csrs_11_V : tlb_1_P1_V;
  wire  _GEN_1026 = 4'h2 == timer[3:0] ? csrs_11_V : tlb_2_P1_V;
  wire  _GEN_1027 = 4'h3 == timer[3:0] ? csrs_11_V : tlb_3_P1_V;
  wire  _GEN_1028 = 4'h4 == timer[3:0] ? csrs_11_V : tlb_4_P1_V;
  wire  _GEN_1029 = 4'h5 == timer[3:0] ? csrs_11_V : tlb_5_P1_V;
  wire  _GEN_1030 = 4'h6 == timer[3:0] ? csrs_11_V : tlb_6_P1_V;
  wire  _GEN_1031 = 4'h7 == timer[3:0] ? csrs_11_V : tlb_7_P1_V;
  wire  _GEN_1032 = 4'h8 == timer[3:0] ? csrs_11_V : tlb_8_P1_V;
  wire  _GEN_1033 = 4'h9 == timer[3:0] ? csrs_11_V : tlb_9_P1_V;
  wire  _GEN_1034 = 4'ha == timer[3:0] ? csrs_11_V : tlb_10_P1_V;
  wire  _GEN_1035 = 4'hb == timer[3:0] ? csrs_11_V : tlb_11_P1_V;
  wire  _GEN_1036 = 4'hc == timer[3:0] ? csrs_11_V : tlb_12_P1_V;
  wire  _GEN_1037 = 4'hd == timer[3:0] ? csrs_11_V : tlb_13_P1_V;
  wire  _GEN_1038 = 4'he == timer[3:0] ? csrs_11_V : tlb_14_P1_V;
  wire  _GEN_1039 = 4'hf == timer[3:0] ? csrs_11_V : tlb_15_P1_V;
  wire  _tlb_0_E_T = ~tlb_0_G;
  wire  _tlb_0_E_T_2 = _tlb_0_E_T & asidMatch_0_1;
  wire  _tlb_0_E_T_5 = _tlb_0_E_T_2 & vaMatch_0_1;
  wire  _tlb_0_E_T_8 = (_tlb_0_E_T | asidMatch_0_1) & vaMatch_0_1;
  wire  _tlb_0_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_0_G | inv_op_decode_2 & _tlb_0_E_T | inv_op_decode_3 &
    _tlb_0_E_T_2 | inv_op_decode_4 & _tlb_0_E_T_5 | inv_op_decode_5 & _tlb_0_E_T_8;
  wire  _tlb_1_E_T = ~tlb_1_G;
  wire  _tlb_1_E_T_2 = _tlb_1_E_T & asidMatch_1_1;
  wire  _tlb_1_E_T_5 = _tlb_1_E_T_2 & vaMatch_1_1;
  wire  _tlb_1_E_T_8 = (_tlb_1_E_T | asidMatch_1_1) & vaMatch_1_1;
  wire  _tlb_1_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_1_G | inv_op_decode_2 & _tlb_1_E_T | inv_op_decode_3 &
    _tlb_1_E_T_2 | inv_op_decode_4 & _tlb_1_E_T_5 | inv_op_decode_5 & _tlb_1_E_T_8;
  wire  _tlb_2_E_T = ~tlb_2_G;
  wire  _tlb_2_E_T_2 = _tlb_2_E_T & asidMatch_2_1;
  wire  _tlb_2_E_T_5 = _tlb_2_E_T_2 & vaMatch_2_1;
  wire  _tlb_2_E_T_8 = (_tlb_2_E_T | asidMatch_2_1) & vaMatch_2_1;
  wire  _tlb_2_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_2_G | inv_op_decode_2 & _tlb_2_E_T | inv_op_decode_3 &
    _tlb_2_E_T_2 | inv_op_decode_4 & _tlb_2_E_T_5 | inv_op_decode_5 & _tlb_2_E_T_8;
  wire  _tlb_3_E_T = ~tlb_3_G;
  wire  _tlb_3_E_T_2 = _tlb_3_E_T & asidMatch_3_1;
  wire  _tlb_3_E_T_5 = _tlb_3_E_T_2 & vaMatch_3_1;
  wire  _tlb_3_E_T_8 = (_tlb_3_E_T | asidMatch_3_1) & vaMatch_3_1;
  wire  _tlb_3_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_3_G | inv_op_decode_2 & _tlb_3_E_T | inv_op_decode_3 &
    _tlb_3_E_T_2 | inv_op_decode_4 & _tlb_3_E_T_5 | inv_op_decode_5 & _tlb_3_E_T_8;
  wire  _tlb_4_E_T = ~tlb_4_G;
  wire  _tlb_4_E_T_2 = _tlb_4_E_T & asidMatch_4_1;
  wire  _tlb_4_E_T_5 = _tlb_4_E_T_2 & vaMatch_4_1;
  wire  _tlb_4_E_T_8 = (_tlb_4_E_T | asidMatch_4_1) & vaMatch_4_1;
  wire  _tlb_4_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_4_G | inv_op_decode_2 & _tlb_4_E_T | inv_op_decode_3 &
    _tlb_4_E_T_2 | inv_op_decode_4 & _tlb_4_E_T_5 | inv_op_decode_5 & _tlb_4_E_T_8;
  wire  _tlb_5_E_T = ~tlb_5_G;
  wire  _tlb_5_E_T_2 = _tlb_5_E_T & asidMatch_5_1;
  wire  _tlb_5_E_T_5 = _tlb_5_E_T_2 & vaMatch_5_1;
  wire  _tlb_5_E_T_8 = (_tlb_5_E_T | asidMatch_5_1) & vaMatch_5_1;
  wire  _tlb_5_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_5_G | inv_op_decode_2 & _tlb_5_E_T | inv_op_decode_3 &
    _tlb_5_E_T_2 | inv_op_decode_4 & _tlb_5_E_T_5 | inv_op_decode_5 & _tlb_5_E_T_8;
  wire  _tlb_6_E_T = ~tlb_6_G;
  wire  _tlb_6_E_T_2 = _tlb_6_E_T & asidMatch_6_1;
  wire  _tlb_6_E_T_5 = _tlb_6_E_T_2 & vaMatch_6_1;
  wire  _tlb_6_E_T_8 = (_tlb_6_E_T | asidMatch_6_1) & vaMatch_6_1;
  wire  _tlb_6_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_6_G | inv_op_decode_2 & _tlb_6_E_T | inv_op_decode_3 &
    _tlb_6_E_T_2 | inv_op_decode_4 & _tlb_6_E_T_5 | inv_op_decode_5 & _tlb_6_E_T_8;
  wire  _tlb_7_E_T = ~tlb_7_G;
  wire  _tlb_7_E_T_2 = _tlb_7_E_T & asidMatch_7_1;
  wire  _tlb_7_E_T_5 = _tlb_7_E_T_2 & vaMatch_7_1;
  wire  _tlb_7_E_T_8 = (_tlb_7_E_T | asidMatch_7_1) & vaMatch_7_1;
  wire  _tlb_7_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_7_G | inv_op_decode_2 & _tlb_7_E_T | inv_op_decode_3 &
    _tlb_7_E_T_2 | inv_op_decode_4 & _tlb_7_E_T_5 | inv_op_decode_5 & _tlb_7_E_T_8;
  wire  _tlb_8_E_T = ~tlb_8_G;
  wire  _tlb_8_E_T_2 = _tlb_8_E_T & asidMatch_8_1;
  wire  _tlb_8_E_T_5 = _tlb_8_E_T_2 & vaMatch_8_1;
  wire  _tlb_8_E_T_8 = (_tlb_8_E_T | asidMatch_8_1) & vaMatch_8_1;
  wire  _tlb_8_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_8_G | inv_op_decode_2 & _tlb_8_E_T | inv_op_decode_3 &
    _tlb_8_E_T_2 | inv_op_decode_4 & _tlb_8_E_T_5 | inv_op_decode_5 & _tlb_8_E_T_8;
  wire  _tlb_9_E_T = ~tlb_9_G;
  wire  _tlb_9_E_T_2 = _tlb_9_E_T & asidMatch_9_1;
  wire  _tlb_9_E_T_5 = _tlb_9_E_T_2 & vaMatch_9_1;
  wire  _tlb_9_E_T_8 = (_tlb_9_E_T | asidMatch_9_1) & vaMatch_9_1;
  wire  _tlb_9_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_9_G | inv_op_decode_2 & _tlb_9_E_T | inv_op_decode_3 &
    _tlb_9_E_T_2 | inv_op_decode_4 & _tlb_9_E_T_5 | inv_op_decode_5 & _tlb_9_E_T_8;
  wire  _tlb_10_E_T = ~tlb_10_G;
  wire  _tlb_10_E_T_2 = _tlb_10_E_T & asidMatch_10_1;
  wire  _tlb_10_E_T_5 = _tlb_10_E_T_2 & vaMatch_10_1;
  wire  _tlb_10_E_T_8 = (_tlb_10_E_T | asidMatch_10_1) & vaMatch_10_1;
  wire  _tlb_10_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_10_G | inv_op_decode_2 & _tlb_10_E_T | inv_op_decode_3
     & _tlb_10_E_T_2 | inv_op_decode_4 & _tlb_10_E_T_5 | inv_op_decode_5 & _tlb_10_E_T_8;
  wire  _tlb_11_E_T = ~tlb_11_G;
  wire  _tlb_11_E_T_2 = _tlb_11_E_T & asidMatch_11_1;
  wire  _tlb_11_E_T_5 = _tlb_11_E_T_2 & vaMatch_11_1;
  wire  _tlb_11_E_T_8 = (_tlb_11_E_T | asidMatch_11_1) & vaMatch_11_1;
  wire  _tlb_11_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_11_G | inv_op_decode_2 & _tlb_11_E_T | inv_op_decode_3
     & _tlb_11_E_T_2 | inv_op_decode_4 & _tlb_11_E_T_5 | inv_op_decode_5 & _tlb_11_E_T_8;
  wire  _tlb_12_E_T = ~tlb_12_G;
  wire  _tlb_12_E_T_2 = _tlb_12_E_T & asidMatch_12_1;
  wire  _tlb_12_E_T_5 = _tlb_12_E_T_2 & vaMatch_12_1;
  wire  _tlb_12_E_T_8 = (_tlb_12_E_T | asidMatch_12_1) & vaMatch_12_1;
  wire  _tlb_12_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_12_G | inv_op_decode_2 & _tlb_12_E_T | inv_op_decode_3
     & _tlb_12_E_T_2 | inv_op_decode_4 & _tlb_12_E_T_5 | inv_op_decode_5 & _tlb_12_E_T_8;
  wire  _tlb_13_E_T = ~tlb_13_G;
  wire  _tlb_13_E_T_2 = _tlb_13_E_T & asidMatch_13_1;
  wire  _tlb_13_E_T_5 = _tlb_13_E_T_2 & vaMatch_13_1;
  wire  _tlb_13_E_T_8 = (_tlb_13_E_T | asidMatch_13_1) & vaMatch_13_1;
  wire  _tlb_13_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_13_G | inv_op_decode_2 & _tlb_13_E_T | inv_op_decode_3
     & _tlb_13_E_T_2 | inv_op_decode_4 & _tlb_13_E_T_5 | inv_op_decode_5 & _tlb_13_E_T_8;
  wire  _tlb_14_E_T = ~tlb_14_G;
  wire  _tlb_14_E_T_2 = _tlb_14_E_T & asidMatch_14_1;
  wire  _tlb_14_E_T_5 = _tlb_14_E_T_2 & vaMatch_14_1;
  wire  _tlb_14_E_T_8 = (_tlb_14_E_T | asidMatch_14_1) & vaMatch_14_1;
  wire  _tlb_14_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_14_G | inv_op_decode_2 & _tlb_14_E_T | inv_op_decode_3
     & _tlb_14_E_T_2 | inv_op_decode_4 & _tlb_14_E_T_5 | inv_op_decode_5 & _tlb_14_E_T_8;
  wire  _tlb_15_E_T = ~tlb_15_G;
  wire  _tlb_15_E_T_2 = _tlb_15_E_T & asidMatch_15_1;
  wire  _tlb_15_E_T_5 = _tlb_15_E_T_2 & vaMatch_15_1;
  wire  _tlb_15_E_T_8 = (_tlb_15_E_T | asidMatch_15_1) & vaMatch_15_1;
  wire  _tlb_15_E_T_19 = inv_op_decode_0 | inv_op_decode_1 & tlb_15_G | inv_op_decode_2 & _tlb_15_E_T | inv_op_decode_3
     & _tlb_15_E_T_2 | inv_op_decode_4 & _tlb_15_E_T_5 | inv_op_decode_5 & _tlb_15_E_T_8;
  wire  _GEN_1040 = 3'h5 == c0_7 ? tlb_0_E & ~_tlb_0_E_T_19 : tlb_0_E;
  wire  _GEN_1041 = 3'h5 == c0_7 ? tlb_1_E & ~_tlb_1_E_T_19 : tlb_1_E;
  wire  _GEN_1042 = 3'h5 == c0_7 ? tlb_2_E & ~_tlb_2_E_T_19 : tlb_2_E;
  wire  _GEN_1043 = 3'h5 == c0_7 ? tlb_3_E & ~_tlb_3_E_T_19 : tlb_3_E;
  wire  _GEN_1044 = 3'h5 == c0_7 ? tlb_4_E & ~_tlb_4_E_T_19 : tlb_4_E;
  wire  _GEN_1045 = 3'h5 == c0_7 ? tlb_5_E & ~_tlb_5_E_T_19 : tlb_5_E;
  wire  _GEN_1046 = 3'h5 == c0_7 ? tlb_6_E & ~_tlb_6_E_T_19 : tlb_6_E;
  wire  _GEN_1047 = 3'h5 == c0_7 ? tlb_7_E & ~_tlb_7_E_T_19 : tlb_7_E;
  wire  _GEN_1048 = 3'h5 == c0_7 ? tlb_8_E & ~_tlb_8_E_T_19 : tlb_8_E;
  wire  _GEN_1049 = 3'h5 == c0_7 ? tlb_9_E & ~_tlb_9_E_T_19 : tlb_9_E;
  wire  _GEN_1050 = 3'h5 == c0_7 ? tlb_10_E & ~_tlb_10_E_T_19 : tlb_10_E;
  wire  _GEN_1051 = 3'h5 == c0_7 ? tlb_11_E & ~_tlb_11_E_T_19 : tlb_11_E;
  wire  _GEN_1052 = 3'h5 == c0_7 ? tlb_12_E & ~_tlb_12_E_T_19 : tlb_12_E;
  wire  _GEN_1053 = 3'h5 == c0_7 ? tlb_13_E & ~_tlb_13_E_T_19 : tlb_13_E;
  wire  _GEN_1054 = 3'h5 == c0_7 ? tlb_14_E & ~_tlb_14_E_T_19 : tlb_14_E;
  wire  _GEN_1055 = 3'h5 == c0_7 ? tlb_15_E & ~_tlb_15_E_T_19 : tlb_15_E;
  wire [18:0] _GEN_1056 = 3'h4 == c0_7 ? _GEN_800 : tlb_0_VPPN;
  wire [18:0] _GEN_1057 = 3'h4 == c0_7 ? _GEN_801 : tlb_1_VPPN;
  wire [18:0] _GEN_1058 = 3'h4 == c0_7 ? _GEN_802 : tlb_2_VPPN;
  wire [18:0] _GEN_1059 = 3'h4 == c0_7 ? _GEN_803 : tlb_3_VPPN;
  wire [18:0] _GEN_1060 = 3'h4 == c0_7 ? _GEN_804 : tlb_4_VPPN;
  wire [18:0] _GEN_1061 = 3'h4 == c0_7 ? _GEN_805 : tlb_5_VPPN;
  wire [18:0] _GEN_1062 = 3'h4 == c0_7 ? _GEN_806 : tlb_6_VPPN;
  wire [18:0] _GEN_1063 = 3'h4 == c0_7 ? _GEN_807 : tlb_7_VPPN;
  wire [18:0] _GEN_1064 = 3'h4 == c0_7 ? _GEN_808 : tlb_8_VPPN;
  wire [18:0] _GEN_1065 = 3'h4 == c0_7 ? _GEN_809 : tlb_9_VPPN;
  wire [18:0] _GEN_1066 = 3'h4 == c0_7 ? _GEN_810 : tlb_10_VPPN;
  wire [18:0] _GEN_1067 = 3'h4 == c0_7 ? _GEN_811 : tlb_11_VPPN;
  wire [18:0] _GEN_1068 = 3'h4 == c0_7 ? _GEN_812 : tlb_12_VPPN;
  wire [18:0] _GEN_1069 = 3'h4 == c0_7 ? _GEN_813 : tlb_13_VPPN;
  wire [18:0] _GEN_1070 = 3'h4 == c0_7 ? _GEN_814 : tlb_14_VPPN;
  wire [18:0] _GEN_1071 = 3'h4 == c0_7 ? _GEN_815 : tlb_15_VPPN;
  wire [5:0] _GEN_1072 = 3'h4 == c0_7 ? _GEN_816 : tlb_0_PS;
  wire [5:0] _GEN_1073 = 3'h4 == c0_7 ? _GEN_817 : tlb_1_PS;
  wire [5:0] _GEN_1074 = 3'h4 == c0_7 ? _GEN_818 : tlb_2_PS;
  wire [5:0] _GEN_1075 = 3'h4 == c0_7 ? _GEN_819 : tlb_3_PS;
  wire [5:0] _GEN_1076 = 3'h4 == c0_7 ? _GEN_820 : tlb_4_PS;
  wire [5:0] _GEN_1077 = 3'h4 == c0_7 ? _GEN_821 : tlb_5_PS;
  wire [5:0] _GEN_1078 = 3'h4 == c0_7 ? _GEN_822 : tlb_6_PS;
  wire [5:0] _GEN_1079 = 3'h4 == c0_7 ? _GEN_823 : tlb_7_PS;
  wire [5:0] _GEN_1080 = 3'h4 == c0_7 ? _GEN_824 : tlb_8_PS;
  wire [5:0] _GEN_1081 = 3'h4 == c0_7 ? _GEN_825 : tlb_9_PS;
  wire [5:0] _GEN_1082 = 3'h4 == c0_7 ? _GEN_826 : tlb_10_PS;
  wire [5:0] _GEN_1083 = 3'h4 == c0_7 ? _GEN_827 : tlb_11_PS;
  wire [5:0] _GEN_1084 = 3'h4 == c0_7 ? _GEN_828 : tlb_12_PS;
  wire [5:0] _GEN_1085 = 3'h4 == c0_7 ? _GEN_829 : tlb_13_PS;
  wire [5:0] _GEN_1086 = 3'h4 == c0_7 ? _GEN_830 : tlb_14_PS;
  wire [5:0] _GEN_1087 = 3'h4 == c0_7 ? _GEN_831 : tlb_15_PS;
  wire  _GEN_1088 = 3'h4 == c0_7 ? _GEN_832 : tlb_0_G;
  wire  _GEN_1089 = 3'h4 == c0_7 ? _GEN_833 : tlb_1_G;
  wire  _GEN_1090 = 3'h4 == c0_7 ? _GEN_834 : tlb_2_G;
  wire  _GEN_1091 = 3'h4 == c0_7 ? _GEN_835 : tlb_3_G;
  wire  _GEN_1092 = 3'h4 == c0_7 ? _GEN_836 : tlb_4_G;
  wire  _GEN_1093 = 3'h4 == c0_7 ? _GEN_837 : tlb_5_G;
  wire  _GEN_1094 = 3'h4 == c0_7 ? _GEN_838 : tlb_6_G;
  wire  _GEN_1095 = 3'h4 == c0_7 ? _GEN_839 : tlb_7_G;
  wire  _GEN_1096 = 3'h4 == c0_7 ? _GEN_840 : tlb_8_G;
  wire  _GEN_1097 = 3'h4 == c0_7 ? _GEN_841 : tlb_9_G;
  wire  _GEN_1098 = 3'h4 == c0_7 ? _GEN_842 : tlb_10_G;
  wire  _GEN_1099 = 3'h4 == c0_7 ? _GEN_843 : tlb_11_G;
  wire  _GEN_1100 = 3'h4 == c0_7 ? _GEN_844 : tlb_12_G;
  wire  _GEN_1101 = 3'h4 == c0_7 ? _GEN_845 : tlb_13_G;
  wire  _GEN_1102 = 3'h4 == c0_7 ? _GEN_846 : tlb_14_G;
  wire  _GEN_1103 = 3'h4 == c0_7 ? _GEN_847 : tlb_15_G;
  wire [9:0] _GEN_1104 = 3'h4 == c0_7 ? _GEN_848 : tlb_0_ASID;
  wire [9:0] _GEN_1105 = 3'h4 == c0_7 ? _GEN_849 : tlb_1_ASID;
  wire [9:0] _GEN_1106 = 3'h4 == c0_7 ? _GEN_850 : tlb_2_ASID;
  wire [9:0] _GEN_1107 = 3'h4 == c0_7 ? _GEN_851 : tlb_3_ASID;
  wire [9:0] _GEN_1108 = 3'h4 == c0_7 ? _GEN_852 : tlb_4_ASID;
  wire [9:0] _GEN_1109 = 3'h4 == c0_7 ? _GEN_853 : tlb_5_ASID;
  wire [9:0] _GEN_1110 = 3'h4 == c0_7 ? _GEN_854 : tlb_6_ASID;
  wire [9:0] _GEN_1111 = 3'h4 == c0_7 ? _GEN_855 : tlb_7_ASID;
  wire [9:0] _GEN_1112 = 3'h4 == c0_7 ? _GEN_856 : tlb_8_ASID;
  wire [9:0] _GEN_1113 = 3'h4 == c0_7 ? _GEN_857 : tlb_9_ASID;
  wire [9:0] _GEN_1114 = 3'h4 == c0_7 ? _GEN_858 : tlb_10_ASID;
  wire [9:0] _GEN_1115 = 3'h4 == c0_7 ? _GEN_859 : tlb_11_ASID;
  wire [9:0] _GEN_1116 = 3'h4 == c0_7 ? _GEN_860 : tlb_12_ASID;
  wire [9:0] _GEN_1117 = 3'h4 == c0_7 ? _GEN_861 : tlb_13_ASID;
  wire [9:0] _GEN_1118 = 3'h4 == c0_7 ? _GEN_862 : tlb_14_ASID;
  wire [9:0] _GEN_1119 = 3'h4 == c0_7 ? _GEN_863 : tlb_15_ASID;
  wire  _GEN_1120 = 3'h4 == c0_7 ? _GEN_864 : _GEN_1040;
  wire  _GEN_1121 = 3'h4 == c0_7 ? _GEN_865 : _GEN_1041;
  wire  _GEN_1122 = 3'h4 == c0_7 ? _GEN_866 : _GEN_1042;
  wire  _GEN_1123 = 3'h4 == c0_7 ? _GEN_867 : _GEN_1043;
  wire  _GEN_1124 = 3'h4 == c0_7 ? _GEN_868 : _GEN_1044;
  wire  _GEN_1125 = 3'h4 == c0_7 ? _GEN_869 : _GEN_1045;
  wire  _GEN_1126 = 3'h4 == c0_7 ? _GEN_870 : _GEN_1046;
  wire  _GEN_1127 = 3'h4 == c0_7 ? _GEN_871 : _GEN_1047;
  wire  _GEN_1128 = 3'h4 == c0_7 ? _GEN_872 : _GEN_1048;
  wire  _GEN_1129 = 3'h4 == c0_7 ? _GEN_873 : _GEN_1049;
  wire  _GEN_1130 = 3'h4 == c0_7 ? _GEN_874 : _GEN_1050;
  wire  _GEN_1131 = 3'h4 == c0_7 ? _GEN_875 : _GEN_1051;
  wire  _GEN_1132 = 3'h4 == c0_7 ? _GEN_876 : _GEN_1052;
  wire  _GEN_1133 = 3'h4 == c0_7 ? _GEN_877 : _GEN_1053;
  wire  _GEN_1134 = 3'h4 == c0_7 ? _GEN_878 : _GEN_1054;
  wire  _GEN_1135 = 3'h4 == c0_7 ? _GEN_879 : _GEN_1055;
  wire [19:0] _GEN_1136 = 3'h4 == c0_7 ? _GEN_880 : tlb_0_P0_PPN;
  wire [19:0] _GEN_1137 = 3'h4 == c0_7 ? _GEN_881 : tlb_1_P0_PPN;
  wire [19:0] _GEN_1138 = 3'h4 == c0_7 ? _GEN_882 : tlb_2_P0_PPN;
  wire [19:0] _GEN_1139 = 3'h4 == c0_7 ? _GEN_883 : tlb_3_P0_PPN;
  wire [19:0] _GEN_1140 = 3'h4 == c0_7 ? _GEN_884 : tlb_4_P0_PPN;
  wire [19:0] _GEN_1141 = 3'h4 == c0_7 ? _GEN_885 : tlb_5_P0_PPN;
  wire [19:0] _GEN_1142 = 3'h4 == c0_7 ? _GEN_886 : tlb_6_P0_PPN;
  wire [19:0] _GEN_1143 = 3'h4 == c0_7 ? _GEN_887 : tlb_7_P0_PPN;
  wire [19:0] _GEN_1144 = 3'h4 == c0_7 ? _GEN_888 : tlb_8_P0_PPN;
  wire [19:0] _GEN_1145 = 3'h4 == c0_7 ? _GEN_889 : tlb_9_P0_PPN;
  wire [19:0] _GEN_1146 = 3'h4 == c0_7 ? _GEN_890 : tlb_10_P0_PPN;
  wire [19:0] _GEN_1147 = 3'h4 == c0_7 ? _GEN_891 : tlb_11_P0_PPN;
  wire [19:0] _GEN_1148 = 3'h4 == c0_7 ? _GEN_892 : tlb_12_P0_PPN;
  wire [19:0] _GEN_1149 = 3'h4 == c0_7 ? _GEN_893 : tlb_13_P0_PPN;
  wire [19:0] _GEN_1150 = 3'h4 == c0_7 ? _GEN_894 : tlb_14_P0_PPN;
  wire [19:0] _GEN_1151 = 3'h4 == c0_7 ? _GEN_895 : tlb_15_P0_PPN;
  wire [1:0] _GEN_1152 = 3'h4 == c0_7 ? _GEN_896 : tlb_0_P0_PLV;
  wire [1:0] _GEN_1153 = 3'h4 == c0_7 ? _GEN_897 : tlb_1_P0_PLV;
  wire [1:0] _GEN_1154 = 3'h4 == c0_7 ? _GEN_898 : tlb_2_P0_PLV;
  wire [1:0] _GEN_1155 = 3'h4 == c0_7 ? _GEN_899 : tlb_3_P0_PLV;
  wire [1:0] _GEN_1156 = 3'h4 == c0_7 ? _GEN_900 : tlb_4_P0_PLV;
  wire [1:0] _GEN_1157 = 3'h4 == c0_7 ? _GEN_901 : tlb_5_P0_PLV;
  wire [1:0] _GEN_1158 = 3'h4 == c0_7 ? _GEN_902 : tlb_6_P0_PLV;
  wire [1:0] _GEN_1159 = 3'h4 == c0_7 ? _GEN_903 : tlb_7_P0_PLV;
  wire [1:0] _GEN_1160 = 3'h4 == c0_7 ? _GEN_904 : tlb_8_P0_PLV;
  wire [1:0] _GEN_1161 = 3'h4 == c0_7 ? _GEN_905 : tlb_9_P0_PLV;
  wire [1:0] _GEN_1162 = 3'h4 == c0_7 ? _GEN_906 : tlb_10_P0_PLV;
  wire [1:0] _GEN_1163 = 3'h4 == c0_7 ? _GEN_907 : tlb_11_P0_PLV;
  wire [1:0] _GEN_1164 = 3'h4 == c0_7 ? _GEN_908 : tlb_12_P0_PLV;
  wire [1:0] _GEN_1165 = 3'h4 == c0_7 ? _GEN_909 : tlb_13_P0_PLV;
  wire [1:0] _GEN_1166 = 3'h4 == c0_7 ? _GEN_910 : tlb_14_P0_PLV;
  wire [1:0] _GEN_1167 = 3'h4 == c0_7 ? _GEN_911 : tlb_15_P0_PLV;
  wire [1:0] _GEN_1168 = 3'h4 == c0_7 ? _GEN_912 : tlb_0_P0_MAT;
  wire [1:0] _GEN_1169 = 3'h4 == c0_7 ? _GEN_913 : tlb_1_P0_MAT;
  wire [1:0] _GEN_1170 = 3'h4 == c0_7 ? _GEN_914 : tlb_2_P0_MAT;
  wire [1:0] _GEN_1171 = 3'h4 == c0_7 ? _GEN_915 : tlb_3_P0_MAT;
  wire [1:0] _GEN_1172 = 3'h4 == c0_7 ? _GEN_916 : tlb_4_P0_MAT;
  wire [1:0] _GEN_1173 = 3'h4 == c0_7 ? _GEN_917 : tlb_5_P0_MAT;
  wire [1:0] _GEN_1174 = 3'h4 == c0_7 ? _GEN_918 : tlb_6_P0_MAT;
  wire [1:0] _GEN_1175 = 3'h4 == c0_7 ? _GEN_919 : tlb_7_P0_MAT;
  wire [1:0] _GEN_1176 = 3'h4 == c0_7 ? _GEN_920 : tlb_8_P0_MAT;
  wire [1:0] _GEN_1177 = 3'h4 == c0_7 ? _GEN_921 : tlb_9_P0_MAT;
  wire [1:0] _GEN_1178 = 3'h4 == c0_7 ? _GEN_922 : tlb_10_P0_MAT;
  wire [1:0] _GEN_1179 = 3'h4 == c0_7 ? _GEN_923 : tlb_11_P0_MAT;
  wire [1:0] _GEN_1180 = 3'h4 == c0_7 ? _GEN_924 : tlb_12_P0_MAT;
  wire [1:0] _GEN_1181 = 3'h4 == c0_7 ? _GEN_925 : tlb_13_P0_MAT;
  wire [1:0] _GEN_1182 = 3'h4 == c0_7 ? _GEN_926 : tlb_14_P0_MAT;
  wire [1:0] _GEN_1183 = 3'h4 == c0_7 ? _GEN_927 : tlb_15_P0_MAT;
  wire  _GEN_1184 = 3'h4 == c0_7 ? _GEN_928 : tlb_0_P0_D;
  wire  _GEN_1185 = 3'h4 == c0_7 ? _GEN_929 : tlb_1_P0_D;
  wire  _GEN_1186 = 3'h4 == c0_7 ? _GEN_930 : tlb_2_P0_D;
  wire  _GEN_1187 = 3'h4 == c0_7 ? _GEN_931 : tlb_3_P0_D;
  wire  _GEN_1188 = 3'h4 == c0_7 ? _GEN_932 : tlb_4_P0_D;
  wire  _GEN_1189 = 3'h4 == c0_7 ? _GEN_933 : tlb_5_P0_D;
  wire  _GEN_1190 = 3'h4 == c0_7 ? _GEN_934 : tlb_6_P0_D;
  wire  _GEN_1191 = 3'h4 == c0_7 ? _GEN_935 : tlb_7_P0_D;
  wire  _GEN_1192 = 3'h4 == c0_7 ? _GEN_936 : tlb_8_P0_D;
  wire  _GEN_1193 = 3'h4 == c0_7 ? _GEN_937 : tlb_9_P0_D;
  wire  _GEN_1194 = 3'h4 == c0_7 ? _GEN_938 : tlb_10_P0_D;
  wire  _GEN_1195 = 3'h4 == c0_7 ? _GEN_939 : tlb_11_P0_D;
  wire  _GEN_1196 = 3'h4 == c0_7 ? _GEN_940 : tlb_12_P0_D;
  wire  _GEN_1197 = 3'h4 == c0_7 ? _GEN_941 : tlb_13_P0_D;
  wire  _GEN_1198 = 3'h4 == c0_7 ? _GEN_942 : tlb_14_P0_D;
  wire  _GEN_1199 = 3'h4 == c0_7 ? _GEN_943 : tlb_15_P0_D;
  wire  _GEN_1200 = 3'h4 == c0_7 ? _GEN_944 : tlb_0_P0_V;
  wire  _GEN_1201 = 3'h4 == c0_7 ? _GEN_945 : tlb_1_P0_V;
  wire  _GEN_1202 = 3'h4 == c0_7 ? _GEN_946 : tlb_2_P0_V;
  wire  _GEN_1203 = 3'h4 == c0_7 ? _GEN_947 : tlb_3_P0_V;
  wire  _GEN_1204 = 3'h4 == c0_7 ? _GEN_948 : tlb_4_P0_V;
  wire  _GEN_1205 = 3'h4 == c0_7 ? _GEN_949 : tlb_5_P0_V;
  wire  _GEN_1206 = 3'h4 == c0_7 ? _GEN_950 : tlb_6_P0_V;
  wire  _GEN_1207 = 3'h4 == c0_7 ? _GEN_951 : tlb_7_P0_V;
  wire  _GEN_1208 = 3'h4 == c0_7 ? _GEN_952 : tlb_8_P0_V;
  wire  _GEN_1209 = 3'h4 == c0_7 ? _GEN_953 : tlb_9_P0_V;
  wire  _GEN_1210 = 3'h4 == c0_7 ? _GEN_954 : tlb_10_P0_V;
  wire  _GEN_1211 = 3'h4 == c0_7 ? _GEN_955 : tlb_11_P0_V;
  wire  _GEN_1212 = 3'h4 == c0_7 ? _GEN_956 : tlb_12_P0_V;
  wire  _GEN_1213 = 3'h4 == c0_7 ? _GEN_957 : tlb_13_P0_V;
  wire  _GEN_1214 = 3'h4 == c0_7 ? _GEN_958 : tlb_14_P0_V;
  wire  _GEN_1215 = 3'h4 == c0_7 ? _GEN_959 : tlb_15_P0_V;
  wire [19:0] _GEN_1216 = 3'h4 == c0_7 ? _GEN_960 : tlb_0_P1_PPN;
  wire [19:0] _GEN_1217 = 3'h4 == c0_7 ? _GEN_961 : tlb_1_P1_PPN;
  wire [19:0] _GEN_1218 = 3'h4 == c0_7 ? _GEN_962 : tlb_2_P1_PPN;
  wire [19:0] _GEN_1219 = 3'h4 == c0_7 ? _GEN_963 : tlb_3_P1_PPN;
  wire [19:0] _GEN_1220 = 3'h4 == c0_7 ? _GEN_964 : tlb_4_P1_PPN;
  wire [19:0] _GEN_1221 = 3'h4 == c0_7 ? _GEN_965 : tlb_5_P1_PPN;
  wire [19:0] _GEN_1222 = 3'h4 == c0_7 ? _GEN_966 : tlb_6_P1_PPN;
  wire [19:0] _GEN_1223 = 3'h4 == c0_7 ? _GEN_967 : tlb_7_P1_PPN;
  wire [19:0] _GEN_1224 = 3'h4 == c0_7 ? _GEN_968 : tlb_8_P1_PPN;
  wire [19:0] _GEN_1225 = 3'h4 == c0_7 ? _GEN_969 : tlb_9_P1_PPN;
  wire [19:0] _GEN_1226 = 3'h4 == c0_7 ? _GEN_970 : tlb_10_P1_PPN;
  wire [19:0] _GEN_1227 = 3'h4 == c0_7 ? _GEN_971 : tlb_11_P1_PPN;
  wire [19:0] _GEN_1228 = 3'h4 == c0_7 ? _GEN_972 : tlb_12_P1_PPN;
  wire [19:0] _GEN_1229 = 3'h4 == c0_7 ? _GEN_973 : tlb_13_P1_PPN;
  wire [19:0] _GEN_1230 = 3'h4 == c0_7 ? _GEN_974 : tlb_14_P1_PPN;
  wire [19:0] _GEN_1231 = 3'h4 == c0_7 ? _GEN_975 : tlb_15_P1_PPN;
  wire [1:0] _GEN_1232 = 3'h4 == c0_7 ? _GEN_976 : tlb_0_P1_PLV;
  wire [1:0] _GEN_1233 = 3'h4 == c0_7 ? _GEN_977 : tlb_1_P1_PLV;
  wire [1:0] _GEN_1234 = 3'h4 == c0_7 ? _GEN_978 : tlb_2_P1_PLV;
  wire [1:0] _GEN_1235 = 3'h4 == c0_7 ? _GEN_979 : tlb_3_P1_PLV;
  wire [1:0] _GEN_1236 = 3'h4 == c0_7 ? _GEN_980 : tlb_4_P1_PLV;
  wire [1:0] _GEN_1237 = 3'h4 == c0_7 ? _GEN_981 : tlb_5_P1_PLV;
  wire [1:0] _GEN_1238 = 3'h4 == c0_7 ? _GEN_982 : tlb_6_P1_PLV;
  wire [1:0] _GEN_1239 = 3'h4 == c0_7 ? _GEN_983 : tlb_7_P1_PLV;
  wire [1:0] _GEN_1240 = 3'h4 == c0_7 ? _GEN_984 : tlb_8_P1_PLV;
  wire [1:0] _GEN_1241 = 3'h4 == c0_7 ? _GEN_985 : tlb_9_P1_PLV;
  wire [1:0] _GEN_1242 = 3'h4 == c0_7 ? _GEN_986 : tlb_10_P1_PLV;
  wire [1:0] _GEN_1243 = 3'h4 == c0_7 ? _GEN_987 : tlb_11_P1_PLV;
  wire [1:0] _GEN_1244 = 3'h4 == c0_7 ? _GEN_988 : tlb_12_P1_PLV;
  wire [1:0] _GEN_1245 = 3'h4 == c0_7 ? _GEN_989 : tlb_13_P1_PLV;
  wire [1:0] _GEN_1246 = 3'h4 == c0_7 ? _GEN_990 : tlb_14_P1_PLV;
  wire [1:0] _GEN_1247 = 3'h4 == c0_7 ? _GEN_991 : tlb_15_P1_PLV;
  wire [1:0] _GEN_1248 = 3'h4 == c0_7 ? _GEN_992 : tlb_0_P1_MAT;
  wire [1:0] _GEN_1249 = 3'h4 == c0_7 ? _GEN_993 : tlb_1_P1_MAT;
  wire [1:0] _GEN_1250 = 3'h4 == c0_7 ? _GEN_994 : tlb_2_P1_MAT;
  wire [1:0] _GEN_1251 = 3'h4 == c0_7 ? _GEN_995 : tlb_3_P1_MAT;
  wire [1:0] _GEN_1252 = 3'h4 == c0_7 ? _GEN_996 : tlb_4_P1_MAT;
  wire [1:0] _GEN_1253 = 3'h4 == c0_7 ? _GEN_997 : tlb_5_P1_MAT;
  wire [1:0] _GEN_1254 = 3'h4 == c0_7 ? _GEN_998 : tlb_6_P1_MAT;
  wire [1:0] _GEN_1255 = 3'h4 == c0_7 ? _GEN_999 : tlb_7_P1_MAT;
  wire [1:0] _GEN_1256 = 3'h4 == c0_7 ? _GEN_1000 : tlb_8_P1_MAT;
  wire [1:0] _GEN_1257 = 3'h4 == c0_7 ? _GEN_1001 : tlb_9_P1_MAT;
  wire [1:0] _GEN_1258 = 3'h4 == c0_7 ? _GEN_1002 : tlb_10_P1_MAT;
  wire [1:0] _GEN_1259 = 3'h4 == c0_7 ? _GEN_1003 : tlb_11_P1_MAT;
  wire [1:0] _GEN_1260 = 3'h4 == c0_7 ? _GEN_1004 : tlb_12_P1_MAT;
  wire [1:0] _GEN_1261 = 3'h4 == c0_7 ? _GEN_1005 : tlb_13_P1_MAT;
  wire [1:0] _GEN_1262 = 3'h4 == c0_7 ? _GEN_1006 : tlb_14_P1_MAT;
  wire [1:0] _GEN_1263 = 3'h4 == c0_7 ? _GEN_1007 : tlb_15_P1_MAT;
  wire  _GEN_1264 = 3'h4 == c0_7 ? _GEN_1008 : tlb_0_P1_D;
  wire  _GEN_1265 = 3'h4 == c0_7 ? _GEN_1009 : tlb_1_P1_D;
  wire  _GEN_1266 = 3'h4 == c0_7 ? _GEN_1010 : tlb_2_P1_D;
  wire  _GEN_1267 = 3'h4 == c0_7 ? _GEN_1011 : tlb_3_P1_D;
  wire  _GEN_1268 = 3'h4 == c0_7 ? _GEN_1012 : tlb_4_P1_D;
  wire  _GEN_1269 = 3'h4 == c0_7 ? _GEN_1013 : tlb_5_P1_D;
  wire  _GEN_1270 = 3'h4 == c0_7 ? _GEN_1014 : tlb_6_P1_D;
  wire  _GEN_1271 = 3'h4 == c0_7 ? _GEN_1015 : tlb_7_P1_D;
  wire  _GEN_1272 = 3'h4 == c0_7 ? _GEN_1016 : tlb_8_P1_D;
  wire  _GEN_1273 = 3'h4 == c0_7 ? _GEN_1017 : tlb_9_P1_D;
  wire  _GEN_1274 = 3'h4 == c0_7 ? _GEN_1018 : tlb_10_P1_D;
  wire  _GEN_1275 = 3'h4 == c0_7 ? _GEN_1019 : tlb_11_P1_D;
  wire  _GEN_1276 = 3'h4 == c0_7 ? _GEN_1020 : tlb_12_P1_D;
  wire  _GEN_1277 = 3'h4 == c0_7 ? _GEN_1021 : tlb_13_P1_D;
  wire  _GEN_1278 = 3'h4 == c0_7 ? _GEN_1022 : tlb_14_P1_D;
  wire  _GEN_1279 = 3'h4 == c0_7 ? _GEN_1023 : tlb_15_P1_D;
  wire  _GEN_1280 = 3'h4 == c0_7 ? _GEN_1024 : tlb_0_P1_V;
  wire  _GEN_1281 = 3'h4 == c0_7 ? _GEN_1025 : tlb_1_P1_V;
  wire  _GEN_1282 = 3'h4 == c0_7 ? _GEN_1026 : tlb_2_P1_V;
  wire  _GEN_1283 = 3'h4 == c0_7 ? _GEN_1027 : tlb_3_P1_V;
  wire  _GEN_1284 = 3'h4 == c0_7 ? _GEN_1028 : tlb_4_P1_V;
  wire  _GEN_1285 = 3'h4 == c0_7 ? _GEN_1029 : tlb_5_P1_V;
  wire  _GEN_1286 = 3'h4 == c0_7 ? _GEN_1030 : tlb_6_P1_V;
  wire  _GEN_1287 = 3'h4 == c0_7 ? _GEN_1031 : tlb_7_P1_V;
  wire  _GEN_1288 = 3'h4 == c0_7 ? _GEN_1032 : tlb_8_P1_V;
  wire  _GEN_1289 = 3'h4 == c0_7 ? _GEN_1033 : tlb_9_P1_V;
  wire  _GEN_1290 = 3'h4 == c0_7 ? _GEN_1034 : tlb_10_P1_V;
  wire  _GEN_1291 = 3'h4 == c0_7 ? _GEN_1035 : tlb_11_P1_V;
  wire  _GEN_1292 = 3'h4 == c0_7 ? _GEN_1036 : tlb_12_P1_V;
  wire  _GEN_1293 = 3'h4 == c0_7 ? _GEN_1037 : tlb_13_P1_V;
  wire  _GEN_1294 = 3'h4 == c0_7 ? _GEN_1038 : tlb_14_P1_V;
  wire  _GEN_1295 = 3'h4 == c0_7 ? _GEN_1039 : tlb_15_P1_V;
  wire  _wbIdx_T_1 = c0_1 == 2'h1;
  wire  _wbIdx_T_2 = c0_1 == 2'h2;
  wire  _wbIdx_T_3 = c0_1 == 2'h3;
  wire [4:0] _wbIdx_T_5 = _wbIdx_T_1 ? 5'h1 : 5'h0;
  wire [4:0] _wbIdx_T_6 = _wbIdx_T_2 ? d : 5'h0;
  wire [4:0] _wbIdx_T_7 = _wbIdx_T_3 ? j : 5'h0;
  wire [4:0] _wbIdx_T_9 = _wbIdx_T_5 | _wbIdx_T_6;
  wire [4:0] wbIdx = _wbIdx_T_9 | _wbIdx_T_7;
  wire  _wbData_T = c0_0 == 3'h0;
  wire  _wbData_T_1 = c0_0 == 3'h1;
  wire  _wbData_T_2 = c0_0 == 3'h2;
  wire  _wbData_T_3 = c0_0 == 3'h3;
  wire  _wbData_T_4 = c0_0 == 3'h4;
  wire  _wbData_T_5 = c0_0 == 3'h5;
  wire  _wbData_T_7 = c0_0 == 3'h6;
  wire  _wbData_T_9 = c0_0 == 3'h7;
  wire [31:0] _wbData_T_10 = _wbData_T ? aluOut : 32'h0;
  wire [31:0] _wbData_T_11 = _wbData_T_1 ? extendData : 32'h0;
  wire [31:0] _wbData_T_12 = _wbData_T_2 ? PC4 : 32'h0;
  wire [31:0] _wbData_T_13 = _wbData_T_3 ? csrRD : 32'h0;
  wire [31:0] _wbData_T_14 = _wbData_T_4 ? csrs_21_TID : 32'h0;
  wire [31:0] _wbData_T_15 = _wbData_T_5 ? timer[63:32] : 32'h0;
  wire [31:0] _wbData_T_16 = _wbData_T_7 ? timer[31:0] : 32'h0;
  wire  _wbData_T_17 = _wbData_T_9 & csrs_25_ROLLB;
  wire [31:0] _wbData_T_18 = _wbData_T_10 | _wbData_T_11;
  wire [31:0] _wbData_T_19 = _wbData_T_18 | _wbData_T_12;
  wire [31:0] _wbData_T_20 = _wbData_T_19 | _wbData_T_13;
  wire [31:0] _wbData_T_21 = _wbData_T_20 | _wbData_T_14;
  wire [31:0] _wbData_T_22 = _wbData_T_21 | _wbData_T_15;
  wire [31:0] _wbData_T_23 = _wbData_T_22 | _wbData_T_16;
  wire [31:0] _GEN_2370 = {{31'd0}, _wbData_T_17};
  wire  _T_1468 = mem_OK & |wbIdx;
  wire  _GEN_2313 = _tlb_E_T | _GEN_248;
  wire  _GEN_2314 = _tlb_E_T ? 1'h0 : _GEN_249;
  wire [1:0] _GEN_2315 = ID_OK & c0_8 ? csrs_1_PPLV : _GEN_251;
  wire  _GEN_2316 = ID_OK & c0_8 ? csrs_1_PIE : _GEN_250;
  wire  _GEN_2319 = ID_OK & c0_8 ? _GEN_2313 : _GEN_248;
  wire  _GEN_2320 = ID_OK & c0_8 ? _GEN_2314 : _GEN_249;
  wire  _GEN_2321 = ID_OK & c0_9 | idle;
  wire [3:0] _ecodeNext_T_1 = ADEF ? 4'h8 : 4'h0;
  wire [1:0] _ecodeNext_T_2 = PIF ? 2'h3 : 2'h0;
  wire [3:0] _ecodeNext_T_3 = INE ? 4'hd : 4'h0;
  wire [3:0] _ecodeNext_T_5 = SYS ? 4'hb : 4'h0;
  wire [3:0] _ecodeNext_T_6 = BRK ? 4'hc : 4'h0;
  wire [3:0] _ecodeNext_T_7 = ALE ? 4'h9 : 4'h0;
  wire [1:0] _ecodeNext_T_10 = PIS ? 2'h2 : 2'h0;
  wire [2:0] _ecodeNext_T_11 = PME ? 3'h4 : 3'h0;
  wire [2:0] _ecodeNext_T_12 = PPI ? 3'h7 : 3'h0;
  wire [5:0] _ecodeNext_T_15 = TLBR ? 6'h3f : 6'h0;
  wire [3:0] _GEN_2371 = {{2'd0}, _ecodeNext_T_2};
  wire [3:0] _ecodeNext_T_17 = _ecodeNext_T_1 | _GEN_2371;
  wire [3:0] _ecodeNext_T_18 = _ecodeNext_T_17 | _ecodeNext_T_3;
  wire [3:0] _ecodeNext_T_20 = _ecodeNext_T_18 | _ecodeNext_T_5;
  wire [3:0] _ecodeNext_T_21 = _ecodeNext_T_20 | _ecodeNext_T_6;
  wire [3:0] _ecodeNext_T_22 = _ecodeNext_T_21 | _ecodeNext_T_7;
  wire [3:0] _GEN_2372 = {{3'd0}, PIL};
  wire [3:0] _ecodeNext_T_24 = _ecodeNext_T_22 | _GEN_2372;
  wire [3:0] _GEN_2373 = {{2'd0}, _ecodeNext_T_10};
  wire [3:0] _ecodeNext_T_25 = _ecodeNext_T_24 | _GEN_2373;
  wire [3:0] _GEN_2374 = {{1'd0}, _ecodeNext_T_11};
  wire [3:0] _ecodeNext_T_26 = _ecodeNext_T_25 | _GEN_2374;
  wire [3:0] _GEN_2375 = {{1'd0}, _ecodeNext_T_12};
  wire [3:0] _ecodeNext_T_27 = _ecodeNext_T_26 | _GEN_2375;
  wire [4:0] _ecodeNext_T_29 = {{1'd0}, _ecodeNext_T_27};
  wire [5:0] _GEN_2376 = {{1'd0}, _ecodeNext_T_29};
  wire [5:0] ecodeNext = _GEN_2376 | _ecodeNext_T_15;
  wire  _T_1477 = _T_1316 & _T_1355;
  wire  _GEN_2330 = TLBR | _GEN_2320;
  wire  _GEN_2340 = _T_1316 & _T_1355 ? _GEN_2330 : _GEN_2320;
  wire  _take_T = rj != rkd;
  wire  _take_T_1 = rj == rkd;
  wire [31:0] _take_T_2 = j == 5'h0 ? 32'h0 : GR_rj_MPORT_data;
  wire [31:0] _take_T_3 = kd == 5'h0 ? 32'h0 : GR_rkd_MPORT_data;
  wire  _take_T_4 = $signed(_take_T_2) >= $signed(_take_T_3);
  wire  _take_T_5 = rj >= rkd;
  wire  _take_T_8 = $signed(_take_T_2) < $signed(_take_T_3);
  wire  _take_T_9 = rj < rkd;
  wire  _GEN_2344 = 3'h2 == brType ? _take_T_1 : 3'h1 == brType & _take_T;
  wire  _GEN_2345 = 3'h3 == brType ? _take_T_4 : _GEN_2344;
  wire  _GEN_2346 = 3'h4 == brType ? _take_T_5 : _GEN_2345;
  wire  _GEN_2347 = 3'h5 == brType ? _take_T_8 : _GEN_2346;
  wire  _GEN_2348 = 3'h6 == brType ? _take_T_9 : _GEN_2347;
  wire [31:0] _PC_T_2 = 3'h7 == brType | _GEN_2348 ? aluOut : PC4;
  wire [31:0] _GEN_2350 = _T_28 ? _PC_T_2 : PC;
  wire [31:0] _GEN_2351 = c0_8 ? csrs_5_PC : _GEN_2350;
  assign GR_rj_MPORT_en = 1'h1;
  assign GR_rj_MPORT_addr = inst[9:5];
  assign GR_rj_MPORT_data = GR[GR_rj_MPORT_addr];
  assign GR_rkd_MPORT_en = 1'h1;
  assign GR_rkd_MPORT_addr = _kd_T_5 ? d : k;
  assign GR_rkd_MPORT_data = GR[GR_rkd_MPORT_addr];
  assign GR_MPORT_data = _wbData_T_23 | _GEN_2370;
  assign GR_MPORT_addr = _wbIdx_T_9 | _wbIdx_T_7;
  assign GR_MPORT_mask = 1'h1;
  assign GR_MPORT_en = _T_1468 & _T_1355;
  assign io_inst_req_valid = reset ? 1'h0 : ~iStallReg & ~dStallReg & IF_OK;
  assign io_inst_req_bits_addr = crmd_DA ? PC : pa;
  assign io_data_req_valid = reset ? 1'h0 : _io_inst_req_valid_T_1 & mem_OK & _EXVA_T & ~preldNop & ~(c0_11 & d[2:0] != 3'h1
    );
  assign io_data_req_bits_wen = _io_data_req_bits_wen_T_4[3:0];
  assign io_data_req_bits_addr = c0_11 & d[4:3] == 2'h2 | ~c0_11 & crmd_PG ? pa_1 : aluOut;
  assign io_data_req_bits_wdata = _io_data_req_bits_wdata_T_2[31:0];
  assign io_data_req_bits_cacop = _T_35 ? 1'h0 : _T_1251;
  assign io_data_req_bits_preld = _T_35 ? 1'h0 : _T_1315;

  assign io_debug_pc = PC;
  assign io_debug_wen = mem_OK & |wbIdx & _T_1355 ? 4'hf : 4'h0;
  assign io_debug_wnum = _wbIdx_T_9 | _wbIdx_T_7;
  assign io_debug_wdata = _wbData_T_23 | _GEN_2370;
  assign io_debug_inst = dStallReg ? inst_reg : io_inst_resp_bits;

  always @(posedge clock) begin
    if (GR_MPORT_en & GR_MPORT_mask) begin
      GR[GR_MPORT_addr] <= GR_MPORT_data;
    end
    if (reset) begin
      idle <= 1'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        idle <= 1'h0;
      end else begin
        idle <= _GEN_2321;
      end
    end else begin
      idle <= _GEN_2321;
    end
    if (reset) begin
      PC <= 32'h1c000000;
    end else if (_T_1477) begin
      if (TLBR) begin
        PC <= _csrRD_T_44;
      end else if (excp) begin
        PC <= _csrRD_T_11;
      end else begin
        PC <= _GEN_2351;
      end
    end
    if (reset) begin
      timer <= 64'h0;
    end else begin
      timer <= _timer_T_1;
    end
    if (reset) begin
      iStallReg <= 1'h0;
    end else begin
      iStallReg <= iStall;
    end
    if (reset) begin
      dStallReg <= 1'h0;
    end else begin
      dStallReg <= dStall;
    end
    if (reset) begin
      crmd_DATM <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T) begin
        crmd_DATM <= _crmd_T_4[8:7];
      end
    end
    if (reset) begin
      crmd_DATF <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T) begin
        crmd_DATF <= _crmd_T_4[6:5];
      end
    end
    if (reset) begin
      crmd_PG <= 1'h0;
    end else if (_T_1316 & _T_1355) begin
      if (TLBR) begin
        crmd_PG <= 1'h0;
      end else begin
        crmd_PG <= _GEN_2319;
      end
    end else begin
      crmd_PG <= _GEN_2319;
    end
    crmd_DA <= reset | _GEN_2340;
    if (reset) begin
      crmd_IE <= 1'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        crmd_IE <= 1'h0;
      end else begin
        crmd_IE <= _GEN_2316;
      end
    end else begin
      crmd_IE <= _GEN_2316;
    end
    if (reset) begin
      crmd_PLV <= 2'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        crmd_PLV <= 2'h0;
      end else begin
        crmd_PLV <= _GEN_2315;
      end
    end else begin
      crmd_PLV <= _GEN_2315;
    end
    if (reset) begin
      csrs_1_PIE <= 1'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        csrs_1_PIE <= crmd_IE;
      end else begin
        csrs_1_PIE <= _GEN_252;
      end
    end else begin
      csrs_1_PIE <= _GEN_252;
    end
    if (reset) begin
      csrs_1_PPLV <= 2'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        csrs_1_PPLV <= crmd_PLV;
      end else begin
        csrs_1_PPLV <= _GEN_253;
      end
    end else begin
      csrs_1_PPLV <= _GEN_253;
    end
    if (reset) begin
      csrs_2_FPE <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_4) begin
        csrs_2_FPE <= _euen_T_3[0];
      end
    end
    if (reset) begin
      csrs_3_LIE <= 13'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_5) begin
        csrs_3_LIE <= _ectl_T_3[12:0];
      end
    end
    if (reset) begin
      csrs_4_Ecode <= 6'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        csrs_4_Ecode <= ecodeNext;
      end
    end
    if (reset) begin
      csrs_4_IS_0 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_6) begin
        if (csrMask[0]) begin
          csrs_4_IS_0 <= rkd[0];
        end
      end
    end
    if (reset) begin
      csrs_4_IS_1 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_6) begin
        if (csrMask[1]) begin
          csrs_4_IS_1 <= rkd[1];
        end
      end
    end
    if (reset) begin
      csrs_4_IS_2 <= 1'h0;
    end else begin
      csrs_4_IS_2 <= io_interrupt[0];
    end
    if (reset) begin
      csrs_4_IS_3 <= 1'h0;
    end else begin
      csrs_4_IS_3 <= io_interrupt[1];
    end
    if (reset) begin
      csrs_4_IS_4 <= 1'h0;
    end else begin
      csrs_4_IS_4 <= io_interrupt[2];
    end
    if (reset) begin
      csrs_4_IS_5 <= 1'h0;
    end else begin
      csrs_4_IS_5 <= io_interrupt[3];
    end
    if (reset) begin
      csrs_4_IS_6 <= 1'h0;
    end else begin
      csrs_4_IS_6 <= io_interrupt[4];
    end
    if (reset) begin
      csrs_4_IS_7 <= 1'h0;
    end else begin
      csrs_4_IS_7 <= io_interrupt[5];
    end
    if (reset) begin
      csrs_4_IS_8 <= 1'h0;
    end else begin
      csrs_4_IS_8 <= io_interrupt[6];
    end
    if (reset) begin
      csrs_4_IS_9 <= 1'h0;
    end else begin
      csrs_4_IS_9 <= io_interrupt[7];
    end
    if (reset) begin
      csrs_4_IS_11 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_40) begin
        if (rkd[0] & csrMask[0]) begin
          csrs_4_IS_11 <= 1'h0;
        end else begin
          csrs_4_IS_11 <= _GEN_228;
        end
      end else begin
        csrs_4_IS_11 <= _GEN_228;
      end
    end else begin
      csrs_4_IS_11 <= _GEN_5;
    end
    if (reset) begin
      csrs_4_IS_12 <= 1'h0;
    end else begin
      csrs_4_IS_12 <= io_ipi;
    end
    if (reset) begin
      csrs_5_PC <= 32'h0;
    end else if (_T_1316 & _T_1355) begin
      if (excp) begin
        csrs_5_PC <= PC;
      end else begin
        csrs_5_PC <= _GEN_258;
      end
    end else begin
      csrs_5_PC <= _GEN_258;
    end
    if (reset) begin
      badv_VAddr <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_9) begin
        badv_VAddr <= _badv_T_3;
      end else begin
        badv_VAddr <= _GEN_176;
      end
    end else begin
      badv_VAddr <= _GEN_176;
    end
    if (reset) begin
      csrs_7_VA <= 26'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_10) begin
        csrs_7_VA <= _eentry_VA_T_3;
      end
    end
    if (reset) begin
      csrs_8_NE <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        if (_miss_T_30) begin
          csrs_8_NE <= 1'h0;
        end else begin
          csrs_8_NE <= 1'h1;
        end
      end else if (3'h2 == c0_7) begin
        csrs_8_NE <= ~_GEN_320;
      end else begin
        csrs_8_NE <= _GEN_261;
      end
    end else begin
      csrs_8_NE <= _GEN_261;
    end
    if (reset) begin
      csrs_8_PS <= 6'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_8_PS <= _GEN_262;
      end else if (3'h2 == c0_7) begin
        csrs_8_PS <= _GEN_545;
      end else begin
        csrs_8_PS <= _GEN_262;
      end
    end else begin
      csrs_8_PS <= _GEN_262;
    end
    if (reset) begin
      csrs_8_Index <= 4'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        if (_miss_T_30) begin
          csrs_8_Index <= _tlbidx_Index_T_34;
        end else begin
          csrs_8_Index <= _GEN_263;
        end
      end else begin
        csrs_8_Index <= _GEN_263;
      end
    end else begin
      csrs_8_Index <= _GEN_263;
    end
    if (reset) begin
      csrs_9_VPPN <= 19'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_9_VPPN <= _GEN_264;
      end else if (3'h2 == c0_7) begin
        csrs_9_VPPN <= _GEN_546;
      end else begin
        csrs_9_VPPN <= _GEN_264;
      end
    end else begin
      csrs_9_VPPN <= _GEN_264;
    end
    if (reset) begin
      csrs_10_PPN <= 24'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_10_PPN <= _GEN_265;
      end else if (3'h2 == c0_7) begin
        csrs_10_PPN <= {{4'd0}, _GEN_547};
      end else begin
        csrs_10_PPN <= _GEN_265;
      end
    end else begin
      csrs_10_PPN <= _GEN_265;
    end
    if (reset) begin
      csrs_10_G <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_10_G <= _GEN_266;
      end else if (3'h2 == c0_7) begin
        csrs_10_G <= _GEN_548;
      end else begin
        csrs_10_G <= _GEN_266;
      end
    end else begin
      csrs_10_G <= _GEN_266;
    end
    if (reset) begin
      csrs_10_MAT <= 2'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_10_MAT <= _GEN_267;
      end else if (3'h2 == c0_7) begin
        csrs_10_MAT <= _GEN_549;
      end else begin
        csrs_10_MAT <= _GEN_267;
      end
    end else begin
      csrs_10_MAT <= _GEN_267;
    end
    if (reset) begin
      csrs_10_PLV <= 2'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_10_PLV <= _GEN_268;
      end else if (3'h2 == c0_7) begin
        csrs_10_PLV <= _GEN_550;
      end else begin
        csrs_10_PLV <= _GEN_268;
      end
    end else begin
      csrs_10_PLV <= _GEN_268;
    end
    if (reset) begin
      csrs_10_D <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_10_D <= _GEN_269;
      end else if (3'h2 == c0_7) begin
        csrs_10_D <= _GEN_551;
      end else begin
        csrs_10_D <= _GEN_269;
      end
    end else begin
      csrs_10_D <= _GEN_269;
    end
    if (reset) begin
      csrs_10_V <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_10_V <= _GEN_270;
      end else if (3'h2 == c0_7) begin
        csrs_10_V <= _GEN_552;
      end else begin
        csrs_10_V <= _GEN_270;
      end
    end else begin
      csrs_10_V <= _GEN_270;
    end
    if (reset) begin
      csrs_11_PPN <= 24'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_11_PPN <= _GEN_271;
      end else if (3'h2 == c0_7) begin
        csrs_11_PPN <= {{4'd0}, _GEN_553};
      end else begin
        csrs_11_PPN <= _GEN_271;
      end
    end else begin
      csrs_11_PPN <= _GEN_271;
    end
    if (reset) begin
      csrs_11_G <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_11_G <= _GEN_272;
      end else if (3'h2 == c0_7) begin
        csrs_11_G <= _GEN_548;
      end else begin
        csrs_11_G <= _GEN_272;
      end
    end else begin
      csrs_11_G <= _GEN_272;
    end
    if (reset) begin
      csrs_11_MAT <= 2'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_11_MAT <= _GEN_273;
      end else if (3'h2 == c0_7) begin
        csrs_11_MAT <= _GEN_555;
      end else begin
        csrs_11_MAT <= _GEN_273;
      end
    end else begin
      csrs_11_MAT <= _GEN_273;
    end
    if (reset) begin
      csrs_11_PLV <= 2'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_11_PLV <= _GEN_274;
      end else if (3'h2 == c0_7) begin
        csrs_11_PLV <= _GEN_556;
      end else begin
        csrs_11_PLV <= _GEN_274;
      end
    end else begin
      csrs_11_PLV <= _GEN_274;
    end
    if (reset) begin
      csrs_11_D <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_11_D <= _GEN_275;
      end else if (3'h2 == c0_7) begin
        csrs_11_D <= _GEN_557;
      end else begin
        csrs_11_D <= _GEN_275;
      end
    end else begin
      csrs_11_D <= _GEN_275;
    end
    if (reset) begin
      csrs_11_V <= 1'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        csrs_11_V <= _GEN_276;
      end else if (3'h2 == c0_7) begin
        csrs_11_V <= _GEN_558;
      end else begin
        csrs_11_V <= _GEN_276;
      end
    end else begin
      csrs_11_V <= _GEN_276;
    end
    if (reset) begin
      asid_ASID <= 10'h0;
    end else if (ID_OK) begin
      if (3'h1 == c0_7) begin
        asid_ASID <= _GEN_277;
      end else if (3'h2 == c0_7) begin
        asid_ASID <= _GEN_559;
      end else begin
        asid_ASID <= _GEN_277;
      end
    end else begin
      asid_ASID <= _GEN_277;
    end
    if (reset) begin
      csrs_13_Base <= 20'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_22) begin
        csrs_13_Base <= _pgdl_Base_T_3;
      end
    end
    if (reset) begin
      csrs_14_Base <= 20'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_24) begin
        csrs_14_Base <= _pgdh_Base_T_3;
      end
    end
    if (reset) begin
      csrs_17_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_32) begin
        csrs_17_Data <= _save0_T_3;
      end
    end
    if (reset) begin
      csrs_18_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_33) begin
        csrs_18_Data <= _save1_T_3;
      end
    end
    if (reset) begin
      csrs_19_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_34) begin
        csrs_19_Data <= _save2_T_3;
      end
    end
    if (reset) begin
      csrs_20_Data <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_35) begin
        csrs_20_Data <= _save3_T_3;
      end
    end
    if (reset) begin
      csrs_21_TID <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_36) begin
        csrs_21_TID <= _tid_T_3;
      end
    end
    if (reset) begin
      csrs_22_InitVal <= 30'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_22_InitVal <= next_InitVal;
      end
    end
    if (reset) begin
      csrs_22_Periodic <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_22_Periodic <= next_Periodic;
      end
    end
    if (reset) begin
      csrs_22_En <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        csrs_22_En <= next_En;
      end
    end
    if (reset) begin
      csrs_23_TimeVal <= 32'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_37) begin
        if (next_En) begin
          csrs_23_TimeVal <= _tval_TimeVal_T_3;
        end else begin
          csrs_23_TimeVal <= _GEN_4;
        end
      end else begin
        csrs_23_TimeVal <= _GEN_4;
      end
    end else begin
      csrs_23_TimeVal <= _GEN_4;
    end
    if (reset) begin
      csrs_25_KLO <= 1'h0;
    end else if (ID_OK & c0_8) begin
      csrs_25_KLO <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_41) begin
        csrs_25_KLO <= _GEN_231;
      end
    end
    if (reset) begin
      csrs_25_ROLLB <= 1'h0;
    end else if (ID_OK & c0_8) begin
      if (~csrs_25_KLO) begin
        csrs_25_ROLLB <= 1'h0;
      end else begin
        csrs_25_ROLLB <= _GEN_291;
      end
    end else begin
      csrs_25_ROLLB <= _GEN_291;
    end
    if (reset) begin
      csrs_26_PA <= 26'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_43) begin
        csrs_26_PA <= _tlbrentry_PA_T_3;
      end
    end
    if (reset) begin
      csrs_27_VSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_VSEG <= _dmw0_VSEG_T_3;
      end
    end
    if (reset) begin
      csrs_27_PSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_PSEG <= _dmw0_PSEG_T_3;
      end
    end
    if (reset) begin
      csrs_27_MAT <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_MAT <= _dmw0_MAT_T_3;
      end
    end
    if (reset) begin
      csrs_27_PLV3 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_PLV3 <= rkd[3] & csrMask[3] | csrs_27_PLV3 & ~csrMask[3];
      end
    end
    if (reset) begin
      csrs_27_PLV0 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_45) begin
        csrs_27_PLV0 <= _T_1415 | csrs_27_PLV0 & ~csrMask[0];
      end
    end
    if (reset) begin
      csrs_28_VSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_VSEG <= _dmw1_VSEG_T_3;
      end
    end
    if (reset) begin
      csrs_28_PSEG <= 3'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_PSEG <= _dmw1_PSEG_T_3;
      end
    end
    if (reset) begin
      csrs_28_MAT <= 2'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_MAT <= _dmw1_MAT_T_3;
      end
    end
    if (reset) begin
      csrs_28_PLV3 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_PLV3 <= rkd[3] & csrMask[3] | csrs_28_PLV3 & ~csrMask[3];
      end
    end
    if (reset) begin
      csrs_28_PLV0 <= 1'h0;
    end else if (ID_OK & c0_4 & |csrMask) begin
      if (_csrRD_T_47) begin
        csrs_28_PLV0 <= _T_1415 | csrs_28_PLV0 & ~csrMask[0];
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_E <= _GEN_624;
          end else begin
            tlb_0_E <= _GEN_1120;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_VPPN <= _GEN_560;
          end else begin
            tlb_0_VPPN <= _GEN_1056;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_PS <= _GEN_576;
          end else begin
            tlb_0_PS <= _GEN_1072;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_G <= _GEN_592;
          end else begin
            tlb_0_G <= _GEN_1088;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_ASID <= _GEN_608;
          end else begin
            tlb_0_ASID <= _GEN_1104;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_E <= _GEN_625;
          end else begin
            tlb_1_E <= _GEN_1121;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_VPPN <= _GEN_561;
          end else begin
            tlb_1_VPPN <= _GEN_1057;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_PS <= _GEN_577;
          end else begin
            tlb_1_PS <= _GEN_1073;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_G <= _GEN_593;
          end else begin
            tlb_1_G <= _GEN_1089;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_ASID <= _GEN_609;
          end else begin
            tlb_1_ASID <= _GEN_1105;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_E <= _GEN_626;
          end else begin
            tlb_2_E <= _GEN_1122;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_VPPN <= _GEN_562;
          end else begin
            tlb_2_VPPN <= _GEN_1058;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_PS <= _GEN_578;
          end else begin
            tlb_2_PS <= _GEN_1074;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_G <= _GEN_594;
          end else begin
            tlb_2_G <= _GEN_1090;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_ASID <= _GEN_610;
          end else begin
            tlb_2_ASID <= _GEN_1106;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_E <= _GEN_627;
          end else begin
            tlb_3_E <= _GEN_1123;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_VPPN <= _GEN_563;
          end else begin
            tlb_3_VPPN <= _GEN_1059;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_PS <= _GEN_579;
          end else begin
            tlb_3_PS <= _GEN_1075;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_G <= _GEN_595;
          end else begin
            tlb_3_G <= _GEN_1091;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_ASID <= _GEN_611;
          end else begin
            tlb_3_ASID <= _GEN_1107;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_E <= _GEN_628;
          end else begin
            tlb_4_E <= _GEN_1124;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_VPPN <= _GEN_564;
          end else begin
            tlb_4_VPPN <= _GEN_1060;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_PS <= _GEN_580;
          end else begin
            tlb_4_PS <= _GEN_1076;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_G <= _GEN_596;
          end else begin
            tlb_4_G <= _GEN_1092;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_ASID <= _GEN_612;
          end else begin
            tlb_4_ASID <= _GEN_1108;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_E <= _GEN_629;
          end else begin
            tlb_5_E <= _GEN_1125;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_VPPN <= _GEN_565;
          end else begin
            tlb_5_VPPN <= _GEN_1061;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_PS <= _GEN_581;
          end else begin
            tlb_5_PS <= _GEN_1077;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_G <= _GEN_597;
          end else begin
            tlb_5_G <= _GEN_1093;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_ASID <= _GEN_613;
          end else begin
            tlb_5_ASID <= _GEN_1109;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_E <= _GEN_630;
          end else begin
            tlb_6_E <= _GEN_1126;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_VPPN <= _GEN_566;
          end else begin
            tlb_6_VPPN <= _GEN_1062;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_PS <= _GEN_582;
          end else begin
            tlb_6_PS <= _GEN_1078;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_G <= _GEN_598;
          end else begin
            tlb_6_G <= _GEN_1094;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_ASID <= _GEN_614;
          end else begin
            tlb_6_ASID <= _GEN_1110;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_E <= _GEN_631;
          end else begin
            tlb_7_E <= _GEN_1127;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_VPPN <= _GEN_567;
          end else begin
            tlb_7_VPPN <= _GEN_1063;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_PS <= _GEN_583;
          end else begin
            tlb_7_PS <= _GEN_1079;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_G <= _GEN_599;
          end else begin
            tlb_7_G <= _GEN_1095;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_ASID <= _GEN_615;
          end else begin
            tlb_7_ASID <= _GEN_1111;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_E <= _GEN_632;
          end else begin
            tlb_8_E <= _GEN_1128;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_VPPN <= _GEN_568;
          end else begin
            tlb_8_VPPN <= _GEN_1064;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_PS <= _GEN_584;
          end else begin
            tlb_8_PS <= _GEN_1080;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_G <= _GEN_600;
          end else begin
            tlb_8_G <= _GEN_1096;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_ASID <= _GEN_616;
          end else begin
            tlb_8_ASID <= _GEN_1112;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_E <= _GEN_633;
          end else begin
            tlb_9_E <= _GEN_1129;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_VPPN <= _GEN_569;
          end else begin
            tlb_9_VPPN <= _GEN_1065;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_PS <= _GEN_585;
          end else begin
            tlb_9_PS <= _GEN_1081;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_G <= _GEN_601;
          end else begin
            tlb_9_G <= _GEN_1097;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_ASID <= _GEN_617;
          end else begin
            tlb_9_ASID <= _GEN_1113;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_E <= _GEN_634;
          end else begin
            tlb_10_E <= _GEN_1130;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_VPPN <= _GEN_570;
          end else begin
            tlb_10_VPPN <= _GEN_1066;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_PS <= _GEN_586;
          end else begin
            tlb_10_PS <= _GEN_1082;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_G <= _GEN_602;
          end else begin
            tlb_10_G <= _GEN_1098;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_ASID <= _GEN_618;
          end else begin
            tlb_10_ASID <= _GEN_1114;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_E <= _GEN_635;
          end else begin
            tlb_11_E <= _GEN_1131;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_VPPN <= _GEN_571;
          end else begin
            tlb_11_VPPN <= _GEN_1067;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_PS <= _GEN_587;
          end else begin
            tlb_11_PS <= _GEN_1083;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_G <= _GEN_603;
          end else begin
            tlb_11_G <= _GEN_1099;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_ASID <= _GEN_619;
          end else begin
            tlb_11_ASID <= _GEN_1115;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_E <= _GEN_636;
          end else begin
            tlb_12_E <= _GEN_1132;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_VPPN <= _GEN_572;
          end else begin
            tlb_12_VPPN <= _GEN_1068;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_PS <= _GEN_588;
          end else begin
            tlb_12_PS <= _GEN_1084;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_G <= _GEN_604;
          end else begin
            tlb_12_G <= _GEN_1100;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_ASID <= _GEN_620;
          end else begin
            tlb_12_ASID <= _GEN_1116;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_E <= _GEN_637;
          end else begin
            tlb_13_E <= _GEN_1133;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_VPPN <= _GEN_573;
          end else begin
            tlb_13_VPPN <= _GEN_1069;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_PS <= _GEN_589;
          end else begin
            tlb_13_PS <= _GEN_1085;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_G <= _GEN_605;
          end else begin
            tlb_13_G <= _GEN_1101;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_ASID <= _GEN_621;
          end else begin
            tlb_13_ASID <= _GEN_1117;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_E <= _GEN_638;
          end else begin
            tlb_14_E <= _GEN_1134;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_VPPN <= _GEN_574;
          end else begin
            tlb_14_VPPN <= _GEN_1070;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_PS <= _GEN_590;
          end else begin
            tlb_14_PS <= _GEN_1086;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_G <= _GEN_606;
          end else begin
            tlb_14_G <= _GEN_1102;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_ASID <= _GEN_622;
          end else begin
            tlb_14_ASID <= _GEN_1118;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_E <= _GEN_639;
          end else begin
            tlb_15_E <= _GEN_1135;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_VPPN <= _GEN_575;
          end else begin
            tlb_15_VPPN <= _GEN_1071;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_PS <= _GEN_591;
          end else begin
            tlb_15_PS <= _GEN_1087;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_G <= _GEN_607;
          end else begin
            tlb_15_G <= _GEN_1103;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_ASID <= _GEN_623;
          end else begin
            tlb_15_ASID <= _GEN_1119;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P1_V <= _GEN_784;
          end else begin
            tlb_0_P1_V <= _GEN_1280;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P1_V <= _GEN_785;
          end else begin
            tlb_1_P1_V <= _GEN_1281;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P1_V <= _GEN_786;
          end else begin
            tlb_2_P1_V <= _GEN_1282;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P1_V <= _GEN_787;
          end else begin
            tlb_3_P1_V <= _GEN_1283;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P1_V <= _GEN_788;
          end else begin
            tlb_4_P1_V <= _GEN_1284;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P1_V <= _GEN_789;
          end else begin
            tlb_5_P1_V <= _GEN_1285;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P1_V <= _GEN_790;
          end else begin
            tlb_6_P1_V <= _GEN_1286;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P1_V <= _GEN_791;
          end else begin
            tlb_7_P1_V <= _GEN_1287;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P1_V <= _GEN_792;
          end else begin
            tlb_8_P1_V <= _GEN_1288;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P1_V <= _GEN_793;
          end else begin
            tlb_9_P1_V <= _GEN_1289;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P1_V <= _GEN_794;
          end else begin
            tlb_10_P1_V <= _GEN_1290;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P1_V <= _GEN_795;
          end else begin
            tlb_11_P1_V <= _GEN_1291;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P1_V <= _GEN_796;
          end else begin
            tlb_12_P1_V <= _GEN_1292;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P1_V <= _GEN_797;
          end else begin
            tlb_13_P1_V <= _GEN_1293;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P1_V <= _GEN_798;
          end else begin
            tlb_14_P1_V <= _GEN_1294;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P1_V <= _GEN_799;
          end else begin
            tlb_15_P1_V <= _GEN_1295;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P0_V <= _GEN_704;
          end else begin
            tlb_0_P0_V <= _GEN_1200;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P0_V <= _GEN_705;
          end else begin
            tlb_1_P0_V <= _GEN_1201;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P0_V <= _GEN_706;
          end else begin
            tlb_2_P0_V <= _GEN_1202;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P0_V <= _GEN_707;
          end else begin
            tlb_3_P0_V <= _GEN_1203;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P0_V <= _GEN_708;
          end else begin
            tlb_4_P0_V <= _GEN_1204;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P0_V <= _GEN_709;
          end else begin
            tlb_5_P0_V <= _GEN_1205;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P0_V <= _GEN_710;
          end else begin
            tlb_6_P0_V <= _GEN_1206;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P0_V <= _GEN_711;
          end else begin
            tlb_7_P0_V <= _GEN_1207;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P0_V <= _GEN_712;
          end else begin
            tlb_8_P0_V <= _GEN_1208;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P0_V <= _GEN_713;
          end else begin
            tlb_9_P0_V <= _GEN_1209;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P0_V <= _GEN_714;
          end else begin
            tlb_10_P0_V <= _GEN_1210;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P0_V <= _GEN_715;
          end else begin
            tlb_11_P0_V <= _GEN_1211;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P0_V <= _GEN_716;
          end else begin
            tlb_12_P0_V <= _GEN_1212;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P0_V <= _GEN_717;
          end else begin
            tlb_13_P0_V <= _GEN_1213;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P0_V <= _GEN_718;
          end else begin
            tlb_14_P0_V <= _GEN_1214;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P0_V <= _GEN_719;
          end else begin
            tlb_15_P0_V <= _GEN_1215;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P1_PLV <= _GEN_736;
          end else begin
            tlb_0_P1_PLV <= _GEN_1232;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P1_PLV <= _GEN_737;
          end else begin
            tlb_1_P1_PLV <= _GEN_1233;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P1_PLV <= _GEN_738;
          end else begin
            tlb_2_P1_PLV <= _GEN_1234;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P1_PLV <= _GEN_739;
          end else begin
            tlb_3_P1_PLV <= _GEN_1235;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P1_PLV <= _GEN_740;
          end else begin
            tlb_4_P1_PLV <= _GEN_1236;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P1_PLV <= _GEN_741;
          end else begin
            tlb_5_P1_PLV <= _GEN_1237;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P1_PLV <= _GEN_742;
          end else begin
            tlb_6_P1_PLV <= _GEN_1238;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P1_PLV <= _GEN_743;
          end else begin
            tlb_7_P1_PLV <= _GEN_1239;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P1_PLV <= _GEN_744;
          end else begin
            tlb_8_P1_PLV <= _GEN_1240;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P1_PLV <= _GEN_745;
          end else begin
            tlb_9_P1_PLV <= _GEN_1241;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P1_PLV <= _GEN_746;
          end else begin
            tlb_10_P1_PLV <= _GEN_1242;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P1_PLV <= _GEN_747;
          end else begin
            tlb_11_P1_PLV <= _GEN_1243;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P1_PLV <= _GEN_748;
          end else begin
            tlb_12_P1_PLV <= _GEN_1244;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P1_PLV <= _GEN_749;
          end else begin
            tlb_13_P1_PLV <= _GEN_1245;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P1_PLV <= _GEN_750;
          end else begin
            tlb_14_P1_PLV <= _GEN_1246;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P1_PLV <= _GEN_751;
          end else begin
            tlb_15_P1_PLV <= _GEN_1247;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P0_PLV <= _GEN_656;
          end else begin
            tlb_0_P0_PLV <= _GEN_1152;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P0_PLV <= _GEN_657;
          end else begin
            tlb_1_P0_PLV <= _GEN_1153;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P0_PLV <= _GEN_658;
          end else begin
            tlb_2_P0_PLV <= _GEN_1154;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P0_PLV <= _GEN_659;
          end else begin
            tlb_3_P0_PLV <= _GEN_1155;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P0_PLV <= _GEN_660;
          end else begin
            tlb_4_P0_PLV <= _GEN_1156;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P0_PLV <= _GEN_661;
          end else begin
            tlb_5_P0_PLV <= _GEN_1157;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P0_PLV <= _GEN_662;
          end else begin
            tlb_6_P0_PLV <= _GEN_1158;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P0_PLV <= _GEN_663;
          end else begin
            tlb_7_P0_PLV <= _GEN_1159;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P0_PLV <= _GEN_664;
          end else begin
            tlb_8_P0_PLV <= _GEN_1160;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P0_PLV <= _GEN_665;
          end else begin
            tlb_9_P0_PLV <= _GEN_1161;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P0_PLV <= _GEN_666;
          end else begin
            tlb_10_P0_PLV <= _GEN_1162;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P0_PLV <= _GEN_667;
          end else begin
            tlb_11_P0_PLV <= _GEN_1163;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P0_PLV <= _GEN_668;
          end else begin
            tlb_12_P0_PLV <= _GEN_1164;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P0_PLV <= _GEN_669;
          end else begin
            tlb_13_P0_PLV <= _GEN_1165;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P0_PLV <= _GEN_670;
          end else begin
            tlb_14_P0_PLV <= _GEN_1166;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P0_PLV <= _GEN_671;
          end else begin
            tlb_15_P0_PLV <= _GEN_1167;
          end
        end
      end
    end
    if (!(dStallReg)) begin
      inst_reg <= io_inst_resp_bits;
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P1_D <= _GEN_768;
          end else begin
            tlb_0_P1_D <= _GEN_1264;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P1_D <= _GEN_769;
          end else begin
            tlb_1_P1_D <= _GEN_1265;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P1_D <= _GEN_770;
          end else begin
            tlb_2_P1_D <= _GEN_1266;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P1_D <= _GEN_771;
          end else begin
            tlb_3_P1_D <= _GEN_1267;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P1_D <= _GEN_772;
          end else begin
            tlb_4_P1_D <= _GEN_1268;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P1_D <= _GEN_773;
          end else begin
            tlb_5_P1_D <= _GEN_1269;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P1_D <= _GEN_774;
          end else begin
            tlb_6_P1_D <= _GEN_1270;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P1_D <= _GEN_775;
          end else begin
            tlb_7_P1_D <= _GEN_1271;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P1_D <= _GEN_776;
          end else begin
            tlb_8_P1_D <= _GEN_1272;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P1_D <= _GEN_777;
          end else begin
            tlb_9_P1_D <= _GEN_1273;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P1_D <= _GEN_778;
          end else begin
            tlb_10_P1_D <= _GEN_1274;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P1_D <= _GEN_779;
          end else begin
            tlb_11_P1_D <= _GEN_1275;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P1_D <= _GEN_780;
          end else begin
            tlb_12_P1_D <= _GEN_1276;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P1_D <= _GEN_781;
          end else begin
            tlb_13_P1_D <= _GEN_1277;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P1_D <= _GEN_782;
          end else begin
            tlb_14_P1_D <= _GEN_1278;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P1_D <= _GEN_783;
          end else begin
            tlb_15_P1_D <= _GEN_1279;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P0_D <= _GEN_688;
          end else begin
            tlb_0_P0_D <= _GEN_1184;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P0_D <= _GEN_689;
          end else begin
            tlb_1_P0_D <= _GEN_1185;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P0_D <= _GEN_690;
          end else begin
            tlb_2_P0_D <= _GEN_1186;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P0_D <= _GEN_691;
          end else begin
            tlb_3_P0_D <= _GEN_1187;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P0_D <= _GEN_692;
          end else begin
            tlb_4_P0_D <= _GEN_1188;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P0_D <= _GEN_693;
          end else begin
            tlb_5_P0_D <= _GEN_1189;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P0_D <= _GEN_694;
          end else begin
            tlb_6_P0_D <= _GEN_1190;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P0_D <= _GEN_695;
          end else begin
            tlb_7_P0_D <= _GEN_1191;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P0_D <= _GEN_696;
          end else begin
            tlb_8_P0_D <= _GEN_1192;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P0_D <= _GEN_697;
          end else begin
            tlb_9_P0_D <= _GEN_1193;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P0_D <= _GEN_698;
          end else begin
            tlb_10_P0_D <= _GEN_1194;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P0_D <= _GEN_699;
          end else begin
            tlb_11_P0_D <= _GEN_1195;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P0_D <= _GEN_700;
          end else begin
            tlb_12_P0_D <= _GEN_1196;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P0_D <= _GEN_701;
          end else begin
            tlb_13_P0_D <= _GEN_1197;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P0_D <= _GEN_702;
          end else begin
            tlb_14_P0_D <= _GEN_1198;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P0_D <= _GEN_703;
          end else begin
            tlb_15_P0_D <= _GEN_1199;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P0_PPN <= _GEN_640;
          end else begin
            tlb_0_P0_PPN <= _GEN_1136;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P0_MAT <= _GEN_672;
          end else begin
            tlb_0_P0_MAT <= _GEN_1168;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P1_PPN <= _GEN_720;
          end else begin
            tlb_0_P1_PPN <= _GEN_1216;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_0_P1_MAT <= _GEN_752;
          end else begin
            tlb_0_P1_MAT <= _GEN_1248;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P0_PPN <= _GEN_641;
          end else begin
            tlb_1_P0_PPN <= _GEN_1137;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P0_MAT <= _GEN_673;
          end else begin
            tlb_1_P0_MAT <= _GEN_1169;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P1_PPN <= _GEN_721;
          end else begin
            tlb_1_P1_PPN <= _GEN_1217;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_1_P1_MAT <= _GEN_753;
          end else begin
            tlb_1_P1_MAT <= _GEN_1249;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P0_PPN <= _GEN_642;
          end else begin
            tlb_2_P0_PPN <= _GEN_1138;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P0_MAT <= _GEN_674;
          end else begin
            tlb_2_P0_MAT <= _GEN_1170;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P1_PPN <= _GEN_722;
          end else begin
            tlb_2_P1_PPN <= _GEN_1218;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_2_P1_MAT <= _GEN_754;
          end else begin
            tlb_2_P1_MAT <= _GEN_1250;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P0_PPN <= _GEN_643;
          end else begin
            tlb_3_P0_PPN <= _GEN_1139;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P0_MAT <= _GEN_675;
          end else begin
            tlb_3_P0_MAT <= _GEN_1171;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P1_PPN <= _GEN_723;
          end else begin
            tlb_3_P1_PPN <= _GEN_1219;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_3_P1_MAT <= _GEN_755;
          end else begin
            tlb_3_P1_MAT <= _GEN_1251;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P0_PPN <= _GEN_644;
          end else begin
            tlb_4_P0_PPN <= _GEN_1140;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P0_MAT <= _GEN_676;
          end else begin
            tlb_4_P0_MAT <= _GEN_1172;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P1_PPN <= _GEN_724;
          end else begin
            tlb_4_P1_PPN <= _GEN_1220;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_4_P1_MAT <= _GEN_756;
          end else begin
            tlb_4_P1_MAT <= _GEN_1252;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P0_PPN <= _GEN_645;
          end else begin
            tlb_5_P0_PPN <= _GEN_1141;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P0_MAT <= _GEN_677;
          end else begin
            tlb_5_P0_MAT <= _GEN_1173;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P1_PPN <= _GEN_725;
          end else begin
            tlb_5_P1_PPN <= _GEN_1221;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_5_P1_MAT <= _GEN_757;
          end else begin
            tlb_5_P1_MAT <= _GEN_1253;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P0_PPN <= _GEN_646;
          end else begin
            tlb_6_P0_PPN <= _GEN_1142;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P0_MAT <= _GEN_678;
          end else begin
            tlb_6_P0_MAT <= _GEN_1174;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P1_PPN <= _GEN_726;
          end else begin
            tlb_6_P1_PPN <= _GEN_1222;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_6_P1_MAT <= _GEN_758;
          end else begin
            tlb_6_P1_MAT <= _GEN_1254;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P0_PPN <= _GEN_647;
          end else begin
            tlb_7_P0_PPN <= _GEN_1143;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P0_MAT <= _GEN_679;
          end else begin
            tlb_7_P0_MAT <= _GEN_1175;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P1_PPN <= _GEN_727;
          end else begin
            tlb_7_P1_PPN <= _GEN_1223;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_7_P1_MAT <= _GEN_759;
          end else begin
            tlb_7_P1_MAT <= _GEN_1255;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P0_PPN <= _GEN_648;
          end else begin
            tlb_8_P0_PPN <= _GEN_1144;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P0_MAT <= _GEN_680;
          end else begin
            tlb_8_P0_MAT <= _GEN_1176;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P1_PPN <= _GEN_728;
          end else begin
            tlb_8_P1_PPN <= _GEN_1224;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_8_P1_MAT <= _GEN_760;
          end else begin
            tlb_8_P1_MAT <= _GEN_1256;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P0_PPN <= _GEN_649;
          end else begin
            tlb_9_P0_PPN <= _GEN_1145;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P0_MAT <= _GEN_681;
          end else begin
            tlb_9_P0_MAT <= _GEN_1177;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P1_PPN <= _GEN_729;
          end else begin
            tlb_9_P1_PPN <= _GEN_1225;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_9_P1_MAT <= _GEN_761;
          end else begin
            tlb_9_P1_MAT <= _GEN_1257;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P0_PPN <= _GEN_650;
          end else begin
            tlb_10_P0_PPN <= _GEN_1146;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P0_MAT <= _GEN_682;
          end else begin
            tlb_10_P0_MAT <= _GEN_1178;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P1_PPN <= _GEN_730;
          end else begin
            tlb_10_P1_PPN <= _GEN_1226;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_10_P1_MAT <= _GEN_762;
          end else begin
            tlb_10_P1_MAT <= _GEN_1258;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P0_PPN <= _GEN_651;
          end else begin
            tlb_11_P0_PPN <= _GEN_1147;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P0_MAT <= _GEN_683;
          end else begin
            tlb_11_P0_MAT <= _GEN_1179;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P1_PPN <= _GEN_731;
          end else begin
            tlb_11_P1_PPN <= _GEN_1227;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_11_P1_MAT <= _GEN_763;
          end else begin
            tlb_11_P1_MAT <= _GEN_1259;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P0_PPN <= _GEN_652;
          end else begin
            tlb_12_P0_PPN <= _GEN_1148;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P0_MAT <= _GEN_684;
          end else begin
            tlb_12_P0_MAT <= _GEN_1180;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P1_PPN <= _GEN_732;
          end else begin
            tlb_12_P1_PPN <= _GEN_1228;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_12_P1_MAT <= _GEN_764;
          end else begin
            tlb_12_P1_MAT <= _GEN_1260;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P0_PPN <= _GEN_653;
          end else begin
            tlb_13_P0_PPN <= _GEN_1149;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P0_MAT <= _GEN_685;
          end else begin
            tlb_13_P0_MAT <= _GEN_1181;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P1_PPN <= _GEN_733;
          end else begin
            tlb_13_P1_PPN <= _GEN_1229;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_13_P1_MAT <= _GEN_765;
          end else begin
            tlb_13_P1_MAT <= _GEN_1261;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P0_PPN <= _GEN_654;
          end else begin
            tlb_14_P0_PPN <= _GEN_1150;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P0_MAT <= _GEN_686;
          end else begin
            tlb_14_P0_MAT <= _GEN_1182;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P1_PPN <= _GEN_734;
          end else begin
            tlb_14_P1_PPN <= _GEN_1230;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_14_P1_MAT <= _GEN_766;
          end else begin
            tlb_14_P1_MAT <= _GEN_1262;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P0_PPN <= _GEN_655;
          end else begin
            tlb_15_P0_PPN <= _GEN_1151;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P0_MAT <= _GEN_687;
          end else begin
            tlb_15_P0_MAT <= _GEN_1183;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P1_PPN <= _GEN_735;
          end else begin
            tlb_15_P1_PPN <= _GEN_1231;
          end
        end
      end
    end
    if (ID_OK) begin
      if (!(3'h1 == c0_7)) begin
        if (!(3'h2 == c0_7)) begin
          if (3'h3 == c0_7) begin
            tlb_15_P1_MAT <= _GEN_767;
          end else begin
            tlb_15_P1_MAT <= _GEN_1263;
          end
        end
      end
    end
  end
endmodule
module SimpleLACoreWrapRAM(
  input         clock,
  input         reset,
  input         io_ipi,
  input  [7:0]  io_interrupt,
  output [31:0] io_debug_pc,
  output [3:0]  io_debug_wen,
  output [4:0]  io_debug_wnum,
  output [31:0] io_debug_wdata,
  output [31:0] io_debug_inst,
  output        io_inst_en,
  output [31:0] io_inst_addr,
  input  [31:0] io_inst_rdata,
  output        io_data_en,
  output [3:0]  io_data_wen,
  output [31:0] io_data_addr,
  output [31:0] io_data_wdata,
  input  [31:0] io_data_rdata
);
  wire  core_clock;
  wire  core_reset;
  wire  core_io_ipi;
  wire [7:0] core_io_interrupt;
  wire  core_io_inst_req_valid;
  wire [31:0] core_io_inst_req_bits_addr;
  wire  core_io_inst_resp_valid;
  wire [31:0] core_io_inst_resp_bits;
  wire  core_io_data_req_valid;
  wire [3:0] core_io_data_req_bits_wen;
  wire [31:0] core_io_data_req_bits_addr;
  wire [31:0] core_io_data_req_bits_wdata;
  wire  core_io_data_req_bits_cacop;
  wire  core_io_data_req_bits_preld;
  wire  core_io_data_resp_valid;
  wire [31:0] core_io_data_resp_bits;
  wire [31:0] core_io_debug_pc;
  wire [3:0] core_io_debug_wen;
  wire [4:0] core_io_debug_wnum;
  wire [31:0] core_io_debug_wdata;
  wire [31:0] core_io_debug_inst;
  SimpleLACore core (
    .clock(core_clock),
    .reset(core_reset),
    .io_ipi(core_io_ipi),
    .io_interrupt(core_io_interrupt),
    .io_inst_req_valid(core_io_inst_req_valid),
    .io_inst_req_bits_addr(core_io_inst_req_bits_addr),
    .io_inst_resp_valid(core_io_inst_resp_valid),
    .io_inst_resp_bits(core_io_inst_resp_bits),
    .io_data_req_valid(core_io_data_req_valid),
    .io_data_req_bits_wen(core_io_data_req_bits_wen),
    .io_data_req_bits_addr(core_io_data_req_bits_addr),
    .io_data_req_bits_wdata(core_io_data_req_bits_wdata),
    .io_data_req_bits_cacop(core_io_data_req_bits_cacop),
    .io_data_req_bits_preld(core_io_data_req_bits_preld),
    .io_data_resp_valid(core_io_data_resp_valid),
    .io_data_resp_bits(core_io_data_resp_bits),
    .io_debug_pc(core_io_debug_pc),
    .io_debug_wen(core_io_debug_wen),
    .io_debug_wnum(core_io_debug_wnum),
    .io_debug_wdata(core_io_debug_wdata),
    .io_debug_inst(core_io_debug_inst)
  );
  assign io_debug_pc = core_io_debug_pc;
  assign io_debug_wen = core_io_debug_wen;
  assign io_debug_wnum = core_io_debug_wnum;
  assign io_debug_wdata = core_io_debug_wdata;
  assign io_debug_inst = core_io_debug_inst;
  assign io_inst_en = core_io_inst_req_valid;
  assign io_inst_addr = core_io_inst_req_bits_addr;
  assign io_data_en = core_io_data_req_valid & ~core_io_data_req_bits_cacop & ~core_io_data_req_bits_preld;
  assign io_data_wen = core_io_data_req_bits_wen;
  assign io_data_addr = core_io_data_req_bits_addr;
  assign io_data_wdata = core_io_data_req_bits_wdata;
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_ipi = io_ipi;
  assign core_io_interrupt = io_interrupt;
  assign core_io_inst_resp_valid = core_io_inst_req_valid;
  assign core_io_inst_resp_bits = io_inst_rdata;
  assign core_io_data_resp_valid = core_io_data_req_valid;
  assign core_io_data_resp_bits = io_data_rdata;
endmodule
